
library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;

entity ctrlrom is
port (addr	:in std_logic_vector (13 downto 0);
        data  :out std_logic_vector (7 downto 0); 
		clk  : in std_logic		);
end ctrlrom;


architecture rtl of ctrlrom is
	type rom_array is array (0 to 16383) of std_logic_vector(7 downto 0);
constant ROM : ROM_ARRAY := (
		x"78",x"A2",x"FF",x"9A",x"A9",x"C9",x"85",x"FB"
		,x"A9",x"F3",x"85",x"FC",x"A9",x"00",x"85",x"FD"
		,x"A9",x"A0",x"85",x"FE",x"A0",x"00",x"A2",x"01"
		,x"CA",x"F0",x"0E",x"B1",x"FB",x"91",x"FD",x"C8"
		,x"D0",x"F9",x"E6",x"FC",x"E6",x"FE",x"4C",x"18"
		,x"C0",x"B1",x"FB",x"91",x"FD",x"C8",x"C0",x"08"
		,x"D0",x"F7",x"20",x"F8",x"E6",x"A9",x"00",x"85"
		,x"02",x"A9",x"B0",x"85",x"03",x"20",x"85",x"E7"
		,x"4C",x"7B",x"C6",x"20",x"21",x"E8",x"AD",x"10"
		,x"B2",x"09",x"24",x"8D",x"10",x"B2",x"29",x"FE"
		,x"8D",x"10",x"B2",x"29",x"FD",x"8D",x"10",x"B2"
		,x"A9",x"3F",x"20",x"BB",x"EC",x"20",x"88",x"C5"
		,x"A9",x"C0",x"20",x"BB",x"EC",x"20",x"88",x"C5"
		,x"A0",x"00",x"20",x"70",x"C0",x"4C",x"81",x"E9"
		,x"20",x"21",x"E8",x"20",x"C6",x"E7",x"A9",x"00"
		,x"A8",x"91",x"02",x"A2",x"00",x"B1",x"02",x"C9"
		,x"08",x"B0",x"64",x"8A",x"20",x"BB",x"EC",x"20"
		,x"10",x"C6",x"A0",x"00",x"B1",x"02",x"20",x"BB"
		,x"EC",x"20",x"4A",x"C6",x"A9",x"00",x"A0",x"01"
		,x"91",x"02",x"C9",x"40",x"B0",x"12",x"A9",x"00"
		,x"20",x"BB",x"EC",x"20",x"A7",x"C5",x"A0",x"01"
		,x"B1",x"02",x"18",x"69",x"01",x"4C",x"98",x"C0"
		,x"A9",x"40",x"20",x"BB",x"EC",x"20",x"10",x"C6"
		,x"A0",x"00",x"B1",x"02",x"20",x"BB",x"EC",x"20"
		,x"4A",x"C6",x"A9",x"00",x"A0",x"01",x"91",x"02"
		,x"C9",x"40",x"B0",x"12",x"A9",x"00",x"20",x"BB"
		,x"EC",x"20",x"A7",x"C5",x"A0",x"01",x"B1",x"02"
		,x"18",x"69",x"01",x"4C",x"C6",x"C0",x"88",x"B1"
		,x"02",x"18",x"69",x"01",x"4C",x"79",x"C0",x"A0"
		,x"02",x"4C",x"7E",x"E9",x"20",x"C6",x"E7",x"A2"
		,x"00",x"A9",x"01",x"20",x"D1",x"EC",x"A0",x"05"
		,x"B1",x"02",x"29",x"07",x"20",x"09",x"ED",x"A0"
		,x"00",x"91",x"02",x"A0",x"04",x"B1",x"02",x"20"
		,x"BB",x"EC",x"20",x"10",x"C6",x"A0",x"03",x"B1"
		,x"02",x"4A",x"4A",x"4A",x"20",x"BB",x"EC",x"20"
		,x"4A",x"C6",x"A0",x"00",x"20",x"00",x"C6",x"A0"
		,x"01",x"91",x"02",x"C8",x"B1",x"02",x"F0",x"0A"
		,x"A0",x"00",x"B1",x"02",x"C8",x"11",x"02",x"4C"
		,x"45",x"C1",x"88",x"AA",x"B1",x"02",x"20",x"D1"
		,x"EC",x"A0",x"02",x"B1",x"02",x"20",x"7C",x"E7"
		,x"20",x"46",x"E7",x"A0",x"01",x"91",x"02",x"A0"
		,x"04",x"B1",x"02",x"20",x"BB",x"EC",x"20",x"10"
		,x"C6",x"A0",x"01",x"B1",x"02",x"20",x"BB",x"EC"
		,x"20",x"A7",x"C5",x"4C",x"82",x"E8",x"20",x"BD"
		,x"E7",x"A2",x"00",x"A9",x"01",x"20",x"D1",x"EC"
		,x"A0",x"05",x"B1",x"02",x"29",x"07",x"20",x"09"
		,x"ED",x"20",x"BB",x"EC",x"AD",x"10",x"B2",x"29"
		,x"FE",x"8D",x"10",x"B2",x"29",x"FD",x"8D",x"10"
		,x"B2",x"A0",x"04",x"B1",x"02",x"4A",x"4A",x"4A"
		,x"20",x"BB",x"EC",x"20",x"4A",x"C6",x"A0",x"05"
		,x"A2",x"00",x"B1",x"02",x"20",x"D1",x"EC",x"A0"
		,x"05",x"B1",x"02",x"20",x"2F",x"E8",x"F0",x"05"
		,x"90",x"03",x"4C",x"87",x"E8",x"A0",x"05",x"B1"
		,x"02",x"20",x"BB",x"EC",x"20",x"10",x"C6",x"A0"
		,x"00",x"20",x"00",x"C6",x"A0",x"01",x"91",x"02"
		,x"C8",x"B1",x"02",x"F0",x"0A",x"A0",x"00",x"B1"
		,x"02",x"C8",x"11",x"02",x"4C",x"DA",x"C1",x"88"
		,x"AA",x"B1",x"02",x"20",x"D1",x"EC",x"A0",x"02"
		,x"B1",x"02",x"20",x"7C",x"E7",x"20",x"46",x"E7"
		,x"A0",x"01",x"91",x"02",x"A0",x"05",x"B1",x"02"
		,x"20",x"BB",x"EC",x"20",x"10",x"C6",x"A0",x"01"
		,x"B1",x"02",x"20",x"BB",x"EC",x"20",x"A7",x"C5"
		,x"A0",x"05",x"B1",x"02",x"18",x"69",x"01",x"91"
		,x"02",x"4C",x"8E",x"C1",x"20",x"E0",x"E7",x"A0"
		,x"05",x"B1",x"02",x"4A",x"4A",x"4A",x"A0",x"03"
		,x"91",x"02",x"C8",x"B1",x"02",x"4A",x"4A",x"4A"
		,x"A0",x"02",x"91",x"02",x"A2",x"00",x"A9",x"FF"
		,x"20",x"D1",x"EC",x"A0",x"07",x"B1",x"02",x"29"
		,x"07",x"20",x"09",x"ED",x"A0",x"01",x"91",x"02"
		,x"A0",x"03",x"A2",x"00",x"B1",x"02",x"20",x"D1"
		,x"EC",x"A0",x"04",x"B1",x"02",x"20",x"2F",x"E8"
		,x"F0",x"05",x"90",x"03",x"4C",x"8C",x"E8",x"A0"
		,x"03",x"A2",x"00",x"B1",x"02",x"20",x"D1",x"EC"
		,x"A0",x"04",x"B1",x"02",x"20",x"2F",x"E8",x"D0"
		,x"26",x"A0",x"01",x"A2",x"00",x"B1",x"02",x"20"
		,x"D1",x"EC",x"A9",x"FF",x"20",x"D1",x"EC",x"A9"
		,x"07",x"20",x"D1",x"EC",x"A0",x"0A",x"B1",x"02"
		,x"29",x"07",x"20",x"36",x"EE",x"20",x"99",x"ED"
		,x"20",x"46",x"E7",x"A0",x"01",x"91",x"02",x"A0"
		,x"06",x"B1",x"02",x"20",x"BB",x"EC",x"20",x"10"
		,x"C6",x"A0",x"03",x"B1",x"02",x"20",x"BB",x"EC"
		,x"20",x"4A",x"C6",x"A0",x"00",x"20",x"00",x"C6"
		,x"A0",x"00",x"91",x"02",x"A0",x"06",x"B1",x"02"
		,x"20",x"BB",x"EC",x"20",x"10",x"C6",x"A0",x"00"
		,x"B1",x"02",x"C8",x"11",x"02",x"20",x"BB",x"EC"
		,x"20",x"A7",x"C5",x"A9",x"FF",x"A0",x"01",x"91"
		,x"02",x"A0",x"03",x"B1",x"02",x"18",x"69",x"01"
		,x"4C",x"26",x"C2",x"20",x"FA",x"E7",x"A2",x"00"
		,x"A0",x"07",x"B1",x"02",x"18",x"A0",x"09",x"71"
		,x"02",x"38",x"E9",x"01",x"A0",x"00",x"91",x"02"
		,x"A0",x"09",x"B1",x"02",x"4A",x"4A",x"4A",x"A0"
		,x"05",x"91",x"02",x"A0",x"00",x"B1",x"02",x"4A"
		,x"4A",x"4A",x"A0",x"04",x"91",x"02",x"A9",x"FF"
		,x"20",x"D1",x"EC",x"A0",x"0B",x"B1",x"02",x"29"
		,x"07",x"20",x"09",x"ED",x"A0",x"03",x"91",x"02"
		,x"A0",x"05",x"A2",x"00",x"B1",x"02",x"20",x"D1"
		,x"EC",x"A0",x"06",x"B1",x"02",x"20",x"2F",x"E8"
		,x"F0",x"05",x"90",x"03",x"4C",x"E4",x"C3",x"A0"
		,x"05",x"A2",x"00",x"B1",x"02",x"20",x"D1",x"EC"
		,x"A0",x"06",x"B1",x"02",x"20",x"2F",x"E8",x"D0"
		,x"26",x"A0",x"03",x"A2",x"00",x"B1",x"02",x"20"
		,x"D1",x"EC",x"A9",x"FF",x"20",x"D1",x"EC",x"A9"
		,x"07",x"20",x"D1",x"EC",x"A0",x"06",x"B1",x"02"
		,x"29",x"07",x"20",x"36",x"EE",x"20",x"99",x"ED"
		,x"20",x"46",x"E7",x"A0",x"03",x"91",x"02",x"AD"
		,x"10",x"B2",x"29",x"FE",x"8D",x"10",x"B2",x"29"
		,x"FD",x"8D",x"10",x"B2",x"A0",x"05",x"B1",x"02"
		,x"20",x"BB",x"EC",x"20",x"4A",x"C6",x"A0",x"0A"
		,x"B1",x"02",x"A0",x"01",x"91",x"02",x"A2",x"00"
		,x"B1",x"02",x"20",x"D1",x"EC",x"A0",x"0A",x"B1"
		,x"02",x"18",x"A0",x"0C",x"71",x"02",x"90",x"01"
		,x"E8",x"20",x"2F",x"E8",x"B0",x"56",x"A0",x"01"
		,x"B1",x"02",x"20",x"BB",x"EC",x"20",x"10",x"C6"
		,x"A0",x"00",x"20",x"00",x"C6",x"A0",x"02",x"91"
		,x"02",x"A0",x"06",x"B1",x"02",x"F0",x"0A",x"A0"
		,x"03",x"B1",x"02",x"88",x"11",x"02",x"4C",x"B5"
		,x"C3",x"A0",x"02",x"AA",x"B1",x"02",x"20",x"D1"
		,x"EC",x"A0",x"05",x"B1",x"02",x"20",x"7C",x"E7"
		,x"20",x"46",x"E7",x"A0",x"02",x"91",x"02",x"88"
		,x"B1",x"02",x"20",x"BB",x"EC",x"20",x"10",x"C6"
		,x"A0",x"02",x"B1",x"02",x"20",x"BB",x"EC",x"20"
		,x"A7",x"C5",x"A0",x"01",x"B1",x"02",x"18",x"69"
		,x"01",x"4C",x"64",x"C3",x"A9",x"FF",x"A0",x"03"
		,x"91",x"02",x"A0",x"05",x"B1",x"02",x"18",x"69"
		,x"01",x"4C",x"F6",x"C2",x"A0",x"0B",x"4C",x"37"
		,x"E7",x"A0",x"02",x"B1",x"02",x"38",x"E9",x"01"
		,x"91",x"02",x"88",x"B1",x"02",x"38",x"E9",x"01"
		,x"91",x"02",x"20",x"E0",x"E7",x"A0",x"08",x"B1"
		,x"02",x"A0",x"03",x"91",x"02",x"A0",x"07",x"B1"
		,x"02",x"A0",x"02",x"91",x"02",x"A0",x"06",x"B1"
		,x"02",x"18",x"A0",x"08",x"71",x"02",x"A0",x"01"
		,x"91",x"02",x"A0",x"04",x"B1",x"02",x"A0",x"00"
		,x"91",x"02",x"20",x"5E",x"C1",x"20",x"E0",x"E7"
		,x"A0",x"08",x"B1",x"02",x"A0",x"03",x"91",x"02"
		,x"A0",x"05",x"B1",x"02",x"18",x"A0",x"07",x"71"
		,x"02",x"A0",x"02",x"91",x"02",x"A0",x"06",x"B1"
		,x"02",x"18",x"A0",x"08",x"71",x"02",x"A0",x"01"
		,x"91",x"02",x"A0",x"04",x"B1",x"02",x"A0",x"00"
		,x"91",x"02",x"20",x"5E",x"C1",x"20",x"D3",x"E7"
		,x"A0",x"07",x"B1",x"02",x"A0",x"02",x"91",x"02"
		,x"A0",x"06",x"B1",x"02",x"A0",x"01",x"91",x"02"
		,x"A0",x"04",x"B1",x"02",x"18",x"A0",x"06",x"71"
		,x"02",x"A0",x"00",x"91",x"02",x"20",x"FC",x"C1"
		,x"20",x"D3",x"E7",x"A0",x"05",x"B1",x"02",x"18"
		,x"A0",x"07",x"71",x"02",x"A0",x"02",x"91",x"02"
		,x"A0",x"06",x"B1",x"02",x"A0",x"01",x"91",x"02"
		,x"A0",x"04",x"B1",x"02",x"18",x"A0",x"06",x"71"
		,x"02",x"A0",x"00",x"91",x"02",x"20",x"FC",x"C1"
		,x"4C",x"82",x"E8",x"A0",x"01",x"B1",x"02",x"8D"
		,x"08",x"A0",x"88",x"B1",x"02",x"8D",x"09",x"A0"
		,x"4C",x"6A",x"E8",x"20",x"E0",x"E7",x"A0",x"05"
		,x"20",x"29",x"E9",x"85",x"06",x"86",x"07",x"18"
		,x"69",x"01",x"90",x"01",x"E8",x"A0",x"04",x"20"
		,x"DB",x"ED",x"A0",x"00",x"B1",x"06",x"A0",x"03"
		,x"91",x"02",x"AA",x"D0",x"03",x"4C",x"87",x"E8"
		,x"B1",x"02",x"C9",x"0A",x"D0",x"11",x"A9",x"08"
		,x"18",x"6D",x"09",x"A0",x"8D",x"09",x"A0",x"A9"
		,x"00",x"8D",x"08",x"A0",x"4C",x"B6",x"C4",x"B1"
		,x"02",x"C9",x"60",x"90",x"0D",x"B1",x"02",x"C9"
		,x"80",x"B0",x"07",x"38",x"B1",x"02",x"E9",x"60"
		,x"91",x"02",x"AD",x"08",x"A0",x"20",x"BB",x"EC"
		,x"20",x"10",x"C6",x"AD",x"09",x"A0",x"4A",x"4A"
		,x"4A",x"20",x"BB",x"EC",x"20",x"4A",x"C6",x"A0"
		,x"03",x"A2",x"00",x"B1",x"02",x"20",x"67",x"E7"
		,x"18",x"69",x"B2",x"A8",x"8A",x"69",x"EF",x"AA"
		,x"98",x"A0",x"00",x"20",x"DB",x"ED",x"A9",x"00"
		,x"A0",x"02",x"91",x"02",x"C9",x"08",x"B0",x"27"
		,x"88",x"20",x"29",x"E9",x"85",x"06",x"86",x"07"
		,x"18",x"69",x"01",x"90",x"01",x"E8",x"A0",x"00"
		,x"20",x"DB",x"ED",x"A0",x"00",x"B1",x"06",x"20"
		,x"BB",x"EC",x"20",x"A7",x"C5",x"A0",x"02",x"B1"
		,x"02",x"18",x"69",x"01",x"4C",x"32",x"C5",x"A9"
		,x"08",x"18",x"6D",x"08",x"A0",x"8D",x"08",x"A0"
		,x"4C",x"B6",x"C4",x"20",x"21",x"E8",x"20",x"BD"
		,x"E7",x"AD",x"10",x"B2",x"09",x"20",x"8D",x"10"
		,x"B2",x"A2",x"00",x"AD",x"10",x"B2",x"29",x"DF"
		,x"8D",x"10",x"B2",x"A0",x"01",x"4C",x"7E",x"E9"
		,x"AD",x"10",x"B2",x"29",x"EF",x"8D",x"10",x"B2"
		,x"29",x"F7",x"8D",x"10",x"B2",x"A9",x"FF",x"8D"
		,x"12",x"B2",x"A0",x"00",x"B1",x"02",x"8D",x"11"
		,x"B2",x"20",x"6B",x"C5",x"4C",x"5B",x"E8",x"AD"
		,x"10",x"B2",x"09",x"10",x"8D",x"10",x"B2",x"29"
		,x"F7",x"8D",x"10",x"B2",x"A9",x"FF",x"8D",x"12"
		,x"B2",x"A0",x"00",x"B1",x"02",x"8D",x"11",x"B2"
		,x"20",x"6B",x"C5",x"4C",x"5B",x"E8",x"20",x"21"
		,x"E8",x"20",x"C6",x"E7",x"A9",x"00",x"8D",x"11"
		,x"B2",x"8D",x"12",x"B2",x"AD",x"10",x"B2",x"09"
		,x"10",x"8D",x"10",x"B2",x"09",x"08",x"8D",x"10"
		,x"B2",x"09",x"20",x"8D",x"10",x"B2",x"EA",x"EA"
		,x"EA",x"AD",x"11",x"B2",x"A0",x"01",x"91",x"02"
		,x"AD",x"10",x"B2",x"29",x"DF",x"8D",x"10",x"B2"
		,x"A2",x"00",x"B1",x"02",x"C8",x"4C",x"7E",x"E9"
		,x"20",x"21",x"E8",x"A0",x"00",x"20",x"C6",x"C5"
		,x"A0",x"00",x"20",x"C6",x"C5",x"4C",x"81",x"E9"
		,x"A0",x"00",x"B1",x"02",x"29",x"7F",x"91",x"02"
		,x"C9",x"40",x"90",x"14",x"38",x"B1",x"02",x"E9"
		,x"40",x"91",x"02",x"AD",x"10",x"B2",x"09",x"01"
		,x"8D",x"10",x"B2",x"29",x"FD",x"4C",x"3A",x"C6"
		,x"AD",x"10",x"B2",x"09",x"02",x"8D",x"10",x"B2"
		,x"29",x"FE",x"8D",x"10",x"B2",x"B1",x"02",x"09"
		,x"40",x"20",x"BB",x"EC",x"20",x"88",x"C5",x"4C"
		,x"5B",x"E8",x"A0",x"00",x"B1",x"02",x"29",x"07"
		,x"91",x"02",x"09",x"B8",x"20",x"BB",x"EC",x"20"
		,x"88",x"C5",x"4C",x"5B",x"E8",x"20",x"21",x"E8"
		,x"20",x"C6",x"E7",x"A0",x"00",x"20",x"F7",x"C8"
		,x"A0",x"00",x"91",x"02",x"20",x"F7",x"C8",x"A0"
		,x"01",x"91",x"02",x"20",x"29",x"E9",x"A0",x"02"
		,x"4C",x"7E",x"E9",x"20",x"21",x"E8",x"A0",x"0B"
		,x"20",x"49",x"EE",x"A0",x"01",x"A9",x"00",x"91"
		,x"02",x"A9",x"02",x"C8",x"91",x"02",x"A0",x"00"
		,x"20",x"E7",x"C8",x"A9",x"D5",x"A2",x"EE",x"20"
		,x"D1",x"EC",x"20",x"1A",x"C9",x"A0",x"00",x"20"
		,x"43",x"C0",x"A9",x"E3",x"A2",x"EE",x"20",x"D1"
		,x"EC",x"20",x"B3",x"C4",x"AD",x"03",x"B2",x"29"
		,x"40",x"F0",x"0D",x"A9",x"00",x"A2",x"EF",x"20"
		,x"D1",x"EC",x"20",x"B3",x"C4",x"4C",x"96",x"C7"
		,x"A9",x"0F",x"A2",x"EF",x"20",x"D1",x"EC",x"20"
		,x"B3",x"C4",x"A9",x"0A",x"A2",x"A0",x"20",x"D1"
		,x"EC",x"A2",x"02",x"A9",x"20",x"20",x"B9",x"E6"
		,x"A9",x"0A",x"A2",x"A0",x"8D",x"40",x"A4",x"8E"
		,x"41",x"A4",x"20",x"ED",x"E7",x"A9",x"2A",x"A2"
		,x"A2",x"A0",x"03",x"91",x"02",x"C8",x"8A",x"91"
		,x"02",x"A9",x"1F",x"A2",x"EF",x"A0",x"01",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"A9",x"01",x"A0"
		,x"00",x"91",x"02",x"20",x"E2",x"C9",x"A0",x"00"
		,x"91",x"02",x"B1",x"02",x"F0",x"3C",x"B1",x"02"
		,x"C9",x"01",x"F0",x"1C",x"C9",x"02",x"F0",x"0B"
		,x"C9",x"03",x"F0",x"07",x"C9",x"0B",x"F0",x"1D"
		,x"4C",x"96",x"C7",x"A9",x"30",x"A2",x"EF",x"20"
		,x"D1",x"EC",x"20",x"B3",x"C4",x"4C",x"96",x"C7"
		,x"A9",x"4D",x"A2",x"EF",x"20",x"D1",x"EC",x"20"
		,x"B3",x"C4",x"4C",x"96",x"C7",x"A9",x"5E",x"A2"
		,x"EF",x"20",x"D1",x"EC",x"20",x"B3",x"C4",x"4C"
		,x"96",x"C7",x"A9",x"72",x"A2",x"EF",x"20",x"D1"
		,x"EC",x"20",x"B3",x"C4",x"20",x"14",x"E8",x"A9"
		,x"2A",x"A2",x"A2",x"A0",x"06",x"91",x"02",x"C8"
		,x"8A",x"91",x"02",x"A9",x"00",x"A0",x"04",x"91"
		,x"02",x"C8",x"A9",x"02",x"91",x"02",x"A9",x"00"
		,x"A0",x"02",x"91",x"02",x"C8",x"A9",x"C0",x"91"
		,x"02",x"A9",x"0B",x"18",x"A6",x"03",x"65",x"02"
		,x"90",x"01",x"E8",x"A0",x"00",x"91",x"02",x"C8"
		,x"8A",x"91",x"02",x"20",x"27",x"CB",x"A0",x"02"
		,x"20",x"29",x"E9",x"20",x"75",x"E7",x"A9",x"87"
		,x"A2",x"EF",x"20",x"D1",x"EC",x"20",x"B3",x"C4"
		,x"A0",x"00",x"20",x"F7",x"C8",x"A0",x"0A",x"91"
		,x"02",x"C9",x"62",x"F0",x"74",x"C9",x"64",x"D0"
		,x"03",x"4C",x"7D",x"C8",x"C9",x"6A",x"D0",x"03"
		,x"4C",x"A6",x"C8",x"C9",x"72",x"D0",x"03",x"4C"
		,x"DA",x"C8",x"C9",x"75",x"D0",x"DA",x"A0",x"00"
		,x"20",x"5D",x"C6",x"A0",x"07",x"20",x"DB",x"ED"
		,x"A0",x"00",x"20",x"5D",x"C6",x"A0",x"05",x"20"
		,x"DB",x"ED",x"A0",x"06",x"20",x"29",x"E9",x"85"
		,x"06",x"86",x"07",x"38",x"E9",x"01",x"B0",x"01"
		,x"CA",x"A0",x"05",x"20",x"DB",x"ED",x"A5",x"06"
		,x"A6",x"07",x"86",x"12",x"05",x"12",x"F0",x"A8"
		,x"A0",x"00",x"20",x"F7",x"C8",x"A0",x"09",x"91"
		,x"02",x"88",x"20",x"29",x"E9",x"85",x"04",x"86"
		,x"05",x"A0",x"09",x"B1",x"02",x"A0",x"00",x"91"
		,x"04",x"A0",x"08",x"20",x"29",x"E9",x"18",x"69"
		,x"01",x"90",x"01",x"E8",x"A0",x"07",x"4C",x"D7"
		,x"C7",x"A0",x"00",x"20",x"5D",x"C6",x"A0",x"07"
		,x"20",x"DB",x"ED",x"A0",x"00",x"20",x"5D",x"C6"
		,x"A0",x"05",x"20",x"DB",x"ED",x"A0",x"06",x"20"
		,x"29",x"E9",x"85",x"06",x"86",x"07",x"38",x"E9"
		,x"01",x"B0",x"01",x"CA",x"A0",x"05",x"20",x"DB"
		,x"ED",x"A5",x"06",x"A6",x"07",x"86",x"12",x"05"
		,x"12",x"D0",x"03",x"4C",x"A0",x"C7",x"A0",x"08"
		,x"20",x"29",x"E9",x"A0",x"00",x"85",x"0A",x"86"
		,x"0B",x"B1",x"0A",x"A0",x"09",x"91",x"02",x"20"
		,x"BB",x"EC",x"20",x"09",x"C9",x"A0",x"08",x"20"
		,x"29",x"E9",x"18",x"69",x"01",x"90",x"01",x"E8"
		,x"A0",x"07",x"4C",x"32",x"C8",x"A0",x"00",x"20"
		,x"5D",x"C6",x"A0",x"07",x"20",x"DB",x"ED",x"20"
		,x"D3",x"E7",x"A0",x"0B",x"20",x"29",x"E9",x"A0"
		,x"01",x"91",x"02",x"C8",x"8A",x"91",x"02",x"A0"
		,x"00",x"20",x"F7",x"C8",x"A0",x"00",x"91",x"02"
		,x"20",x"48",x"C9",x"4C",x"A0",x"C7",x"A0",x"00"
		,x"20",x"5D",x"C6",x"A0",x"07",x"20",x"DB",x"ED"
		,x"20",x"D3",x"E7",x"A9",x"0A",x"18",x"A6",x"03"
		,x"65",x"02",x"90",x"01",x"E8",x"A0",x"01",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"98",x"A0",x"00"
		,x"91",x"02",x"20",x"48",x"C9",x"A0",x"08",x"20"
		,x"29",x"E9",x"A0",x"01",x"20",x"DB",x"ED",x"20"
		,x"75",x"E7",x"A9",x"92",x"A2",x"EF",x"20",x"D1"
		,x"EC",x"20",x"1A",x"C9",x"4C",x"A0",x"C7",x"20"
		,x"21",x"E8",x"A2",x"01",x"A9",x"0F",x"8D",x"04"
		,x"B1",x"8E",x"05",x"B1",x"4C",x"81",x"E9",x"20"
		,x"21",x"E8",x"AD",x"02",x"B1",x"29",x"01",x"F0"
		,x"F9",x"A2",x"00",x"AD",x"00",x"B1",x"4C",x"81"
		,x"E9",x"AD",x"02",x"B1",x"29",x"02",x"F0",x"F9"
		,x"A0",x"00",x"B1",x"02",x"8D",x"00",x"B1",x"4C"
		,x"5B",x"E8",x"20",x"BD",x"E7",x"A0",x"02",x"20"
		,x"29",x"E9",x"85",x"06",x"86",x"07",x"18",x"69"
		,x"01",x"90",x"01",x"E8",x"A0",x"01",x"20",x"DB"
		,x"ED",x"A0",x"00",x"B1",x"06",x"91",x"02",x"AA"
		,x"D0",x"03",x"4C",x"78",x"E8",x"B1",x"02",x"20"
		,x"BB",x"EC",x"20",x"09",x"C9",x"4C",x"1D",x"C9"
		,x"A9",x"00",x"20",x"BB",x"EC",x"20",x"D3",x"E7"
		,x"A0",x"04",x"B1",x"02",x"48",x"38",x"E9",x"01"
		,x"91",x"02",x"68",x"AA",x"D0",x"03",x"4C",x"8C"
		,x"E8",x"20",x"E0",x"E7",x"A0",x"0A",x"20",x"29"
		,x"E9",x"85",x"06",x"86",x"07",x"18",x"69",x"01"
		,x"90",x"01",x"E8",x"A0",x"09",x"20",x"DB",x"ED"
		,x"A0",x"00",x"B1",x"06",x"A0",x"02",x"91",x"02"
		,x"C8",x"A9",x"00",x"91",x"02",x"A9",x"04",x"18"
		,x"A6",x"03",x"65",x"02",x"90",x"01",x"E8",x"A0"
		,x"00",x"91",x"02",x"C8",x"8A",x"91",x"02",x"A2"
		,x"00",x"A9",x"10",x"20",x"CD",x"E5",x"A0",x"01"
		,x"B1",x"02",x"D0",x"0A",x"A9",x"9B",x"A2",x"EF"
		,x"20",x"D1",x"EC",x"20",x"1A",x"C9",x"A5",x"02"
		,x"A6",x"03",x"20",x"D1",x"EC",x"20",x"1A",x"C9"
		,x"A9",x"9D",x"A2",x"EF",x"20",x"D1",x"EC",x"20"
		,x"1A",x"C9",x"A0",x"03",x"18",x"A9",x"01",x"71"
		,x"02",x"91",x"02",x"C9",x"10",x"D0",x"81",x"A9"
		,x"9F",x"A2",x"EF",x"20",x"D1",x"EC",x"20",x"1A"
		,x"C9",x"A9",x"00",x"A0",x"03",x"91",x"02",x"4C"
		,x"50",x"C9",x"A0",x"1D",x"20",x"49",x"EE",x"AD"
		,x"40",x"A4",x"AE",x"41",x"A4",x"20",x"D1",x"EC"
		,x"A0",x"00",x"20",x"DE",x"DD",x"A0",x"1E",x"91"
		,x"02",x"C9",x"00",x"F0",x"07",x"A2",x"00",x"B1"
		,x"02",x"4C",x"22",x"CB",x"20",x"14",x"E8",x"A9"
		,x"16",x"18",x"A6",x"03",x"65",x"02",x"90",x"01"
		,x"E8",x"A0",x"06",x"91",x"02",x"C8",x"8A",x"91"
		,x"02",x"A9",x"0A",x"18",x"A6",x"03",x"65",x"02"
		,x"90",x"01",x"E8",x"A0",x"04",x"91",x"02",x"C8"
		,x"8A",x"91",x"02",x"A0",x"29",x"20",x"29",x"E9"
		,x"A0",x"02",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A9",x"24",x"18",x"A6",x"03",x"65",x"02",x"90"
		,x"01",x"E8",x"A0",x"00",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"20",x"28",x"DB",x"A0",x"1E",x"91"
		,x"02",x"B1",x"02",x"F0",x"07",x"A2",x"00",x"B1"
		,x"02",x"4C",x"22",x"CB",x"A0",x"1C",x"B1",x"02"
		,x"C8",x"11",x"02",x"F0",x"15",x"20",x"29",x"E9"
		,x"18",x"69",x"0B",x"90",x"01",x"E8",x"A0",x"00"
		,x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"29",x"10"
		,x"F0",x"07",x"A2",x"00",x"A9",x"02",x"4C",x"22"
		,x"CB",x"A0",x"23",x"20",x"29",x"E9",x"85",x"04"
		,x"86",x"05",x"A0",x"1F",x"B1",x"02",x"29",x"01"
		,x"A0",x"14",x"91",x"04",x"A0",x"25",x"20",x"E9"
		,x"EC",x"A0",x"1F",x"20",x"29",x"E9",x"18",x"69"
		,x"14",x"90",x"01",x"E8",x"A0",x"01",x"20",x"1C"
		,x"E9",x"86",x"05",x"85",x"04",x"A9",x"00",x"AA"
		,x"20",x"28",x"EA",x"A0",x"23",x"20",x"29",x"E9"
		,x"18",x"69",x"1A",x"90",x"01",x"E8",x"A0",x"01"
		,x"20",x"1C",x"E9",x"A0",x"00",x"84",x"04",x"84"
		,x"05",x"20",x"04",x"EA",x"A0",x"08",x"20",x"E4"
		,x"ED",x"A0",x"25",x"20",x"E9",x"EC",x"A0",x"1F"
		,x"20",x"29",x"E9",x"18",x"69",x"1C",x"90",x"01"
		,x"E8",x"A0",x"03",x"20",x"32",x"E9",x"A0",x"04"
		,x"20",x"E4",x"ED",x"A0",x"25",x"20",x"E9",x"EC"
		,x"A2",x"00",x"86",x"04",x"86",x"05",x"8A",x"A8"
		,x"20",x"E4",x"ED",x"A0",x"23",x"20",x"29",x"E9"
		,x"85",x"04",x"86",x"05",x"A9",x"01",x"A0",x"15"
		,x"91",x"04",x"A8",x"20",x"29",x"E9",x"85",x"04"
		,x"86",x"05",x"A0",x"01",x"85",x"0A",x"86",x"0B"
		,x"B1",x"0A",x"18",x"69",x"01",x"91",x"04",x"A2"
		,x"00",x"8A",x"A0",x"24",x"4C",x"37",x"E7",x"A0"
		,x"0F",x"20",x"49",x"EE",x"A0",x"16",x"20",x"E9"
		,x"EC",x"AD",x"40",x"A4",x"AE",x"41",x"A4",x"20"
		,x"D1",x"EC",x"A0",x"14",x"20",x"29",x"E9",x"85"
		,x"04",x"86",x"05",x"A9",x"00",x"A8",x"91",x"04"
		,x"C8",x"91",x"04",x"B1",x"02",x"88",x"11",x"02"
		,x"D0",x"06",x"AA",x"A9",x"0A",x"4C",x"FD",x"CE"
		,x"20",x"63",x"DF",x"29",x"01",x"D0",x"10",x"A0"
		,x"01",x"20",x"29",x"E9",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"B1",x"0A",x"AA",x"D0",x"07",x"A2"
		,x"00",x"A9",x"01",x"4C",x"FD",x"CE",x"A0",x"1A"
		,x"20",x"29",x"E9",x"A0",x"14",x"85",x"0A",x"86"
		,x"0B",x"B1",x"0A",x"29",x"80",x"F0",x"03",x"4C"
		,x"F9",x"CE",x"A0",x"1A",x"20",x"29",x"E9",x"A0"
		,x"14",x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"29"
		,x"01",x"D0",x"06",x"AA",x"A9",x"05",x"4C",x"FD"
		,x"CE",x"A0",x"1A",x"20",x"29",x"E9",x"A0",x"07"
		,x"20",x"32",x"E9",x"20",x"28",x"EA",x"A0",x"1E"
		,x"20",x"29",x"E9",x"A0",x"03",x"20",x"32",x"E9"
		,x"20",x"AF",x"EB",x"A0",x"07",x"20",x"0C",x"EE"
		,x"A0",x"18",x"20",x"E9",x"EC",x"A0",x"0C",x"20"
		,x"49",x"E9",x"20",x"56",x"EE",x"20",x"59",x"EC"
		,x"F0",x"0A",x"A0",x"08",x"20",x"29",x"E9",x"A0"
		,x"15",x"20",x"DB",x"ED",x"A0",x"16",x"B1",x"02"
		,x"88",x"11",x"02",x"D0",x"03",x"4C",x"E4",x"CE"
		,x"A0",x"1A",x"20",x"29",x"E9",x"A0",x"03",x"20"
		,x"32",x"E9",x"20",x"28",x"EA",x"A2",x"01",x"A9"
		,x"00",x"85",x"04",x"85",x"05",x"A9",x"FF",x"20"
		,x"B0",x"E8",x"20",x"28",x"EA",x"A2",x"00",x"86"
		,x"04",x"86",x"05",x"8A",x"20",x"91",x"E9",x"D0"
		,x"03",x"4C",x"F2",x"CD",x"A0",x"1A",x"20",x"29"
		,x"E9",x"85",x"0A",x"86",x"0B",x"A0",x"15",x"B1"
		,x"0A",x"38",x"E9",x"01",x"91",x"0A",x"AA",x"F0"
		,x"17",x"A0",x"1A",x"20",x"29",x"E9",x"A0",x"13"
		,x"20",x"32",x"E9",x"A0",x"01",x"20",x"97",x"E9"
		,x"A0",x"0B",x"20",x"0C",x"EE",x"4C",x"E5",x"CC"
		,x"A0",x"1A",x"20",x"29",x"E9",x"A0",x"03",x"20"
		,x"32",x"E9",x"20",x"28",x"EA",x"A2",x"00",x"86"
		,x"04",x"86",x"05",x"8A",x"20",x"91",x"E9",x"F0"
		,x"0D",x"A0",x"1A",x"20",x"29",x"E9",x"A0",x"0B"
		,x"20",x"32",x"E9",x"4C",x"76",x"CC",x"A0",x"1A"
		,x"20",x"29",x"E9",x"A0",x"0F",x"20",x"32",x"E9"
		,x"20",x"28",x"EA",x"20",x"6B",x"D4",x"A0",x"0F"
		,x"20",x"0C",x"EE",x"A0",x"12",x"20",x"49",x"E9"
		,x"C9",x"02",x"8A",x"E9",x"00",x"A5",x"04",x"E9"
		,x"00",x"A5",x"05",x"E9",x"00",x"B0",x"03",x"4C"
		,x"E8",x"CE",x"A0",x"12",x"20",x"49",x"E9",x"20"
		,x"28",x"EA",x"A0",x"05",x"20",x"29",x"E9",x"A0"
		,x"0F",x"20",x"32",x"E9",x"20",x"53",x"EC",x"F0"
		,x"03",x"4C",x"E8",x"CE",x"A0",x"1C",x"20",x"E9"
		,x"EC",x"A0",x"14",x"20",x"49",x"E9",x"A0",x"0C"
		,x"20",x"E4",x"ED",x"A0",x"12",x"20",x"49",x"E9"
		,x"20",x"28",x"EA",x"20",x"97",x"D6",x"A0",x"0B"
		,x"20",x"0C",x"EE",x"A0",x"1A",x"20",x"29",x"E9"
		,x"85",x"04",x"86",x"05",x"A0",x"01",x"20",x"29"
		,x"E9",x"A0",x"02",x"85",x"0A",x"86",x"0B",x"B1"
		,x"0A",x"A0",x"15",x"91",x"04",x"A0",x"1C",x"20"
		,x"E9",x"EC",x"A0",x"10",x"20",x"49",x"E9",x"A0"
		,x"10",x"20",x"E4",x"ED",x"A0",x"16",x"20",x"29"
		,x"E9",x"8A",x"4A",x"A0",x"04",x"91",x"02",x"B1"
		,x"02",x"D0",x"03",x"4C",x"C2",x"CD",x"A2",x"00"
		,x"B1",x"02",x"20",x"D1",x"EC",x"A0",x"1C",x"20"
		,x"29",x"E9",x"A0",x"15",x"85",x"0A",x"86",x"0B"
		,x"A2",x"00",x"B1",x"0A",x"20",x"2F",x"E8",x"90"
		,x"13",x"F0",x"11",x"A0",x"1A",x"20",x"29",x"E9"
		,x"A0",x"15",x"85",x"0A",x"86",x"0B",x"B1",x"0A"
		,x"A0",x"04",x"91",x"02",x"20",x"07",x"E8",x"A0"
		,x"0A",x"20",x"29",x"E9",x"A0",x"05",x"91",x"02"
		,x"C8",x"8A",x"91",x"02",x"A0",x"15",x"20",x"49"
		,x"E9",x"A0",x"01",x"20",x"0C",x"EE",x"A0",x"0B"
		,x"B1",x"02",x"A0",x"00",x"91",x"02",x"20",x"69"
		,x"DF",x"C9",x"00",x"F0",x"03",x"4C",x"E8",x"CE"
		,x"A0",x"1A",x"20",x"29",x"E9",x"20",x"D1",x"EC"
		,x"A0",x"15",x"85",x"0A",x"86",x"0B",x"A2",x"00"
		,x"B1",x"0A",x"20",x"D1",x"EC",x"A0",x"08",x"B1"
		,x"02",x"38",x"E9",x"01",x"B0",x"01",x"CA",x"20"
		,x"36",x"EE",x"A0",x"15",x"20",x"C3",x"ED",x"A0"
		,x"1A",x"20",x"29",x"E9",x"20",x"D1",x"EC",x"A0"
		,x"13",x"20",x"32",x"E9",x"20",x"28",x"EA",x"A0"
		,x"0A",x"A2",x"00",x"B1",x"02",x"38",x"E9",x"01"
		,x"B0",x"01",x"CA",x"A0",x"00",x"84",x"04",x"84"
		,x"05",x"20",x"91",x"E8",x"A0",x"10",x"20",x"E4"
		,x"ED",x"A0",x"04",x"B1",x"02",x"AA",x"A9",x"00"
		,x"20",x"54",x"E7",x"C8",x"20",x"DB",x"ED",x"4C"
		,x"75",x"CE",x"20",x"07",x"E8",x"A0",x"21",x"20"
		,x"29",x"E9",x"18",x"69",x"16",x"90",x"01",x"E8"
		,x"A0",x"05",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A0",x"15",x"20",x"49",x"E9",x"A0",x"01",x"20"
		,x"0C",x"EE",x"A9",x"01",x"A0",x"00",x"91",x"02"
		,x"20",x"69",x"DF",x"C9",x"00",x"F0",x"03",x"4C"
		,x"E8",x"CE",x"A2",x"02",x"A9",x"00",x"20",x"D1"
		,x"EC",x"A0",x"1C",x"20",x"29",x"E9",x"A0",x"01"
		,x"20",x"1C",x"E9",x"A8",x"8A",x"29",x"01",x"AA"
		,x"98",x"20",x"36",x"EE",x"A0",x"05",x"20",x"DB"
		,x"ED",x"20",x"D1",x"EC",x"A0",x"18",x"20",x"29"
		,x"E9",x"20",x"2F",x"E8",x"90",x"0C",x"F0",x"0A"
		,x"A0",x"16",x"20",x"29",x"E9",x"A0",x"05",x"20"
		,x"DB",x"ED",x"20",x"E0",x"E7",x"A0",x"07",x"20"
		,x"29",x"E9",x"A0",x"02",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"A0",x"1E",x"20",x"29",x"E9",x"18"
		,x"69",x"16",x"90",x"01",x"E8",x"20",x"D1",x"EC"
		,x"A0",x"20",x"20",x"29",x"E9",x"A0",x"03",x"20"
		,x"32",x"E9",x"20",x"28",x"EA",x"A2",x"01",x"A9"
		,x"00",x"85",x"04",x"85",x"05",x"A9",x"FF",x"20"
		,x"B0",x"E8",x"20",x"1E",x"E7",x"A0",x"00",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"A0",x"0A",x"20"
		,x"29",x"E9",x"20",x"7F",x"E6",x"A0",x"05",x"B1"
		,x"02",x"A0",x"02",x"18",x"71",x"02",x"91",x"02"
		,x"A0",x"06",x"B1",x"02",x"A0",x"03",x"71",x"02"
		,x"91",x"02",x"A0",x"1A",x"20",x"29",x"E9",x"20"
		,x"D1",x"EC",x"A0",x"03",x"20",x"32",x"E9",x"20"
		,x"28",x"EA",x"A0",x"0C",x"20",x"29",x"E9",x"A0"
		,x"00",x"84",x"04",x"84",x"05",x"20",x"91",x"E8"
		,x"A0",x"00",x"20",x"E4",x"ED",x"A0",x"14",x"20"
		,x"29",x"E9",x"85",x"04",x"86",x"05",x"A0",x"01"
		,x"20",x"1C",x"E9",x"85",x"0A",x"86",x"0B",x"A0"
		,x"06",x"20",x"29",x"E9",x"18",x"65",x"0A",x"85"
		,x"0A",x"8A",x"65",x"0B",x"AA",x"A5",x"0A",x"A0"
		,x"00",x"91",x"04",x"C8",x"8A",x"91",x"04",x"A0"
		,x"06",x"20",x"29",x"E9",x"A0",x"15",x"20",x"21"
		,x"EE",x"4C",x"DC",x"CB",x"AA",x"4C",x"FD",x"CE"
		,x"A0",x"1A",x"20",x"29",x"E9",x"85",x"0A",x"86"
		,x"0B",x"A0",x"14",x"B1",x"0A",x"09",x"80",x"91"
		,x"0A",x"A2",x"00",x"A9",x"07",x"A0",x"1B",x"4C"
		,x"37",x"E7",x"20",x"BD",x"E7",x"A9",x"00",x"A8"
		,x"91",x"02",x"B1",x"02",x"D0",x"26",x"A0",x"02"
		,x"20",x"29",x"E9",x"85",x"04",x"86",x"05",x"A9"
		,x"00",x"A0",x"14",x"91",x"04",x"AD",x"40",x"A4"
		,x"AE",x"41",x"A4",x"85",x"04",x"86",x"05",x"A0"
		,x"01",x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"38"
		,x"E9",x"01",x"91",x"04",x"A0",x"00",x"A2",x"00"
		,x"B1",x"02",x"4C",x"78",x"E8",x"20",x"ED",x"E7"
		,x"AD",x"40",x"A4",x"AE",x"41",x"A4",x"20",x"D1"
		,x"EC",x"A0",x"01",x"B1",x"02",x"88",x"11",x"02"
		,x"D0",x"06",x"AA",x"A9",x"0A",x"4C",x"67",x"D1"
		,x"20",x"63",x"DF",x"29",x"01",x"D0",x"10",x"A0"
		,x"01",x"20",x"29",x"E9",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"B1",x"0A",x"AA",x"D0",x"07",x"A2"
		,x"00",x"A9",x"01",x"4C",x"67",x"D1",x"A0",x"0C"
		,x"20",x"29",x"E9",x"A0",x"14",x"85",x"0A",x"86"
		,x"0B",x"B1",x"0A",x"29",x"80",x"F0",x"03",x"4C"
		,x"63",x"D1",x"A0",x"0A",x"20",x"49",x"E9",x"20"
		,x"28",x"EA",x"A0",x"10",x"20",x"29",x"E9",x"A0"
		,x"07",x"20",x"32",x"E9",x"20",x"59",x"EC",x"F0"
		,x"0F",x"A0",x"0C",x"20",x"29",x"E9",x"A0",x"07"
		,x"20",x"32",x"E9",x"A0",x"07",x"20",x"0C",x"EE"
		,x"A0",x"0E",x"20",x"E9",x"EC",x"A0",x"0C",x"20"
		,x"49",x"E9",x"A0",x"00",x"20",x"E4",x"ED",x"A0"
		,x"0C",x"20",x"29",x"E9",x"85",x"04",x"86",x"05"
		,x"A9",x"01",x"A0",x"15",x"91",x"04",x"A0",x"0A"
		,x"20",x"49",x"E9",x"D0",x"03",x"4C",x"4C",x"D1"
		,x"A0",x"0A",x"20",x"49",x"E9",x"A0",x"01",x"20"
		,x"5A",x"E9",x"20",x"28",x"EA",x"A2",x"00",x"86"
		,x"04",x"86",x"05",x"A9",x"09",x"20",x"17",x"EB"
		,x"A0",x"07",x"20",x"0C",x"EE",x"A0",x"01",x"20"
		,x"29",x"E9",x"A0",x"02",x"85",x"0A",x"86",x"0B"
		,x"B1",x"0A",x"91",x"02",x"A0",x"0E",x"20",x"E9"
		,x"EC",x"A0",x"04",x"A2",x"00",x"B1",x"02",x"20"
		,x"D1",x"EC",x"A0",x"0B",x"B1",x"02",x"20",x"D1"
		,x"EC",x"A0",x"08",x"B1",x"02",x"20",x"C6",x"EE"
		,x"20",x"36",x"EE",x"A0",x"15",x"20",x"C3",x"ED"
		,x"A0",x"0A",x"20",x"49",x"E9",x"20",x"28",x"EA"
		,x"A0",x"06",x"A2",x"00",x"B1",x"02",x"A0",x"00"
		,x"86",x"04",x"86",x"05",x"20",x"DF",x"EB",x"A0"
		,x"07",x"20",x"0C",x"EE",x"A0",x"0C",x"20",x"29"
		,x"E9",x"A0",x"0B",x"20",x"32",x"E9",x"A0",x"03"
		,x"20",x"0C",x"EE",x"A0",x"0A",x"20",x"49",x"E9"
		,x"20",x"40",x"EA",x"A0",x"01",x"20",x"5A",x"E9"
		,x"A0",x"07",x"20",x"0C",x"EE",x"20",x"4F",x"EA"
		,x"20",x"D0",x"EB",x"F0",x"0E",x"A0",x"06",x"20"
		,x"49",x"E9",x"20",x"28",x"EA",x"20",x"6B",x"D4"
		,x"4C",x"4E",x"D0",x"A0",x"06",x"20",x"49",x"E9"
		,x"C9",x"02",x"8A",x"E9",x"00",x"A5",x"04",x"E9"
		,x"00",x"A5",x"05",x"E9",x"00",x"B0",x"03",x"4C"
		,x"52",x"D1",x"A0",x"06",x"20",x"49",x"E9",x"20"
		,x"28",x"EA",x"A0",x"05",x"20",x"29",x"E9",x"A0"
		,x"0F",x"20",x"32",x"E9",x"20",x"53",x"EC",x"F0"
		,x"03",x"4C",x"52",x"D1",x"A0",x"0E",x"20",x"E9"
		,x"EC",x"A0",x"08",x"20",x"49",x"E9",x"A0",x"0C"
		,x"20",x"E4",x"ED",x"A0",x"0E",x"20",x"E9",x"EC"
		,x"A0",x"08",x"20",x"49",x"E9",x"20",x"28",x"EA"
		,x"20",x"97",x"D6",x"20",x"28",x"EA",x"A0",x"08"
		,x"A2",x"00",x"B1",x"02",x"A0",x"00",x"86",x"04"
		,x"86",x"05",x"20",x"91",x"E8",x"20",x"28",x"EA"
		,x"A0",x"12",x"20",x"29",x"E9",x"A0",x"15",x"85"
		,x"0A",x"86",x"0B",x"A2",x"00",x"B1",x"0A",x"86"
		,x"04",x"86",x"05",x"20",x"AF",x"EB",x"A0",x"10"
		,x"20",x"E4",x"ED",x"A0",x"0C",x"20",x"29",x"E9"
		,x"A0",x"03",x"20",x"32",x"E9",x"20",x"28",x"EA"
		,x"A2",x"01",x"A9",x"00",x"85",x"04",x"85",x"05"
		,x"A9",x"FF",x"20",x"B0",x"E8",x"20",x"D0",x"EB"
		,x"F0",x"32",x"20",x"07",x"E8",x"A0",x"13",x"20"
		,x"29",x"E9",x"18",x"69",x"16",x"90",x"01",x"E8"
		,x"A0",x"05",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A0",x"13",x"20",x"29",x"E9",x"A0",x"13",x"20"
		,x"32",x"E9",x"A0",x"01",x"20",x"0C",x"EE",x"A9"
		,x"01",x"A0",x"00",x"91",x"02",x"20",x"69",x"DF"
		,x"C9",x"00",x"D0",x"06",x"A2",x"00",x"8A",x"4C"
		,x"67",x"D1",x"A0",x"0C",x"20",x"29",x"E9",x"85"
		,x"0A",x"86",x"0B",x"A0",x"14",x"B1",x"0A",x"09"
		,x"80",x"91",x"0A",x"A2",x"00",x"A9",x"07",x"A0"
		,x"0D",x"4C",x"37",x"E7",x"A0",x"0D",x"20",x"49"
		,x"EE",x"AD",x"40",x"A4",x"AE",x"41",x"A4",x"20"
		,x"D1",x"EC",x"A0",x"01",x"B1",x"02",x"88",x"11"
		,x"02",x"D0",x"06",x"AA",x"A9",x"0A",x"4C",x"E7"
		,x"D3",x"A0",x"03",x"20",x"E9",x"EC",x"A2",x"02"
		,x"A9",x"20",x"20",x"B9",x"E6",x"20",x"3A",x"DE"
		,x"29",x"01",x"F0",x"07",x"A2",x"00",x"A9",x"01"
		,x"4C",x"E7",x"D3",x"AA",x"85",x"04",x"85",x"05"
		,x"A0",x"0A",x"20",x"0C",x"EE",x"20",x"28",x"EA"
		,x"20",x"FE",x"D6",x"A0",x"0E",x"91",x"02",x"B1"
		,x"02",x"D0",x"35",x"A0",x"01",x"20",x"29",x"E9"
		,x"E8",x"A0",x"E2",x"85",x"0A",x"86",x"0B",x"B1"
		,x"0A",x"F0",x"25",x"A0",x"01",x"20",x"29",x"E9"
		,x"18",x"69",x"E6",x"90",x"01",x"E8",x"E8",x"A0"
		,x"03",x"20",x"32",x"E9",x"A0",x"0A",x"20",x"0C"
		,x"EE",x"A0",x"0D",x"20",x"49",x"E9",x"20",x"28"
		,x"EA",x"20",x"FE",x"D6",x"A0",x"0E",x"91",x"02"
		,x"A0",x"0E",x"B1",x"02",x"D0",x"06",x"AA",x"A9"
		,x"0B",x"4C",x"E7",x"D3",x"A0",x"01",x"20",x"29"
		,x"E9",x"85",x"04",x"86",x"05",x"A0",x"0E",x"B1"
		,x"02",x"A0",x"00",x"91",x"04",x"A0",x"03",x"20"
		,x"E9",x"EC",x"A0",x"10",x"B1",x"02",x"C9",x"03"
		,x"D0",x"12",x"A8",x"20",x"29",x"E9",x"18",x"69"
		,x"44",x"90",x"01",x"E8",x"A0",x"03",x"20",x"32"
		,x"E9",x"4C",x"42",x"D2",x"A0",x"03",x"20",x"29"
		,x"E9",x"18",x"69",x"36",x"90",x"01",x"E8",x"A0"
		,x"01",x"20",x"1C",x"E9",x"A0",x"00",x"84",x"04"
		,x"84",x"05",x"A0",x"08",x"20",x"E4",x"ED",x"A0"
		,x"01",x"20",x"29",x"E9",x"85",x"04",x"86",x"05"
		,x"A0",x"01",x"20",x"29",x"E9",x"A0",x"2D",x"85"
		,x"0A",x"86",x"0B",x"B1",x"0A",x"A0",x"02",x"91"
		,x"04",x"88",x"20",x"29",x"E9",x"85",x"04",x"86"
		,x"05",x"A0",x"01",x"20",x"29",x"E9",x"A0",x"30"
		,x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"A0",x"03"
		,x"91",x"04",x"A0",x"03",x"20",x"E9",x"EC",x"A0"
		,x"0F",x"20",x"49",x"E9",x"20",x"28",x"EA",x"A0"
		,x"07",x"20",x"29",x"E9",x"18",x"69",x"2E",x"90"
		,x"01",x"E8",x"A0",x"01",x"20",x"1C",x"E9",x"A0"
		,x"00",x"84",x"04",x"84",x"05",x"20",x"91",x"E8"
		,x"A0",x"10",x"20",x"E4",x"ED",x"A0",x"01",x"20"
		,x"29",x"E9",x"85",x"04",x"86",x"05",x"A0",x"01"
		,x"20",x"29",x"E9",x"18",x"69",x"31",x"90",x"01"
		,x"E8",x"A0",x"01",x"20",x"1C",x"E9",x"A0",x"04"
		,x"91",x"04",x"C8",x"8A",x"91",x"04",x"A0",x"01"
		,x"20",x"29",x"E9",x"A0",x"0B",x"20",x"32",x"E9"
		,x"20",x"28",x"EA",x"A0",x"05",x"20",x"29",x"E9"
		,x"A0",x"03",x"85",x"0A",x"86",x"0B",x"A2",x"00"
		,x"B1",x"0A",x"86",x"04",x"86",x"05",x"20",x"A8"
		,x"E9",x"20",x"28",x"EA",x"A0",x"05",x"20",x"29"
		,x"E9",x"A0",x"13",x"20",x"32",x"E9",x"20",x"91"
		,x"E8",x"A0",x"06",x"20",x"0C",x"EE",x"A0",x"0E"
		,x"B1",x"02",x"C9",x"03",x"D0",x"26",x"A8",x"20"
		,x"E9",x"EC",x"A0",x"03",x"20",x"29",x"E9",x"18"
		,x"69",x"4C",x"90",x"01",x"E8",x"A0",x"03",x"20"
		,x"32",x"E9",x"A0",x"14",x"20",x"E4",x"ED",x"A0"
		,x"03",x"20",x"E9",x"EC",x"A0",x"0B",x"20",x"49"
		,x"E9",x"4C",x"5B",x"D3",x"A0",x"03",x"20",x"E9"
		,x"EC",x"A0",x"0B",x"20",x"49",x"E9",x"A0",x"14"
		,x"20",x"E4",x"ED",x"A0",x"03",x"20",x"E9",x"EC"
		,x"A0",x"03",x"20",x"29",x"E9",x"A0",x"05",x"20"
		,x"1C",x"E9",x"20",x"45",x"ED",x"20",x"D1",x"EC"
		,x"A0",x"0D",x"20",x"49",x"E9",x"20",x"56",x"EE"
		,x"20",x"91",x"E8",x"A0",x"18",x"20",x"E4",x"ED"
		,x"A0",x"01",x"20",x"29",x"E9",x"18",x"69",x"40"
		,x"90",x"01",x"E8",x"A0",x"03",x"20",x"32",x"E9"
		,x"A0",x"02",x"20",x"0C",x"EE",x"A0",x"05",x"20"
		,x"49",x"E9",x"20",x"CE",x"E8",x"F0",x"1B",x"A0"
		,x"01",x"20",x"29",x"E9",x"18",x"69",x"33",x"90"
		,x"01",x"E8",x"A0",x"01",x"20",x"1C",x"E9",x"A0"
		,x"00",x"84",x"04",x"84",x"05",x"A0",x"02",x"20"
		,x"0C",x"EE",x"A0",x"03",x"20",x"E9",x"EC",x"A0"
		,x"07",x"20",x"49",x"E9",x"20",x"28",x"EA",x"A0"
		,x"07",x"20",x"29",x"E9",x"A0",x"1B",x"20",x"32"
		,x"E9",x"20",x"AF",x"EB",x"20",x"28",x"EA",x"A0"
		,x"13",x"20",x"49",x"E9",x"20",x"91",x"E8",x"20"
		,x"28",x"EA",x"A0",x"07",x"20",x"29",x"E9",x"A0"
		,x"02",x"85",x"0A",x"86",x"0B",x"A2",x"00",x"B1"
		,x"0A",x"A0",x"00",x"86",x"04",x"86",x"05",x"20"
		,x"DF",x"EB",x"A0",x"02",x"20",x"97",x"E9",x"A0"
		,x"0C",x"20",x"E4",x"ED",x"A2",x"00",x"8A",x"A0"
		,x"0F",x"4C",x"37",x"E7",x"20",x"E0",x"E7",x"AD"
		,x"40",x"A4",x"AE",x"41",x"A4",x"20",x"D1",x"EC"
		,x"A0",x"01",x"20",x"29",x"E9",x"A0",x"1F",x"20"
		,x"32",x"E9",x"A0",x"02",x"20",x"0C",x"EE",x"A0"
		,x"05",x"20",x"49",x"E9",x"20",x"28",x"EA",x"A0"
		,x"0D",x"20",x"49",x"E9",x"20",x"FE",x"E9",x"F0"
		,x"49",x"A0",x"09",x"20",x"49",x"E9",x"F0",x"42"
		,x"20",x"07",x"E8",x"A0",x"08",x"20",x"29",x"E9"
		,x"18",x"69",x"20",x"90",x"01",x"E8",x"A0",x"05"
		,x"91",x"02",x"C8",x"8A",x"91",x"02",x"A0",x"10"
		,x"20",x"49",x"E9",x"A0",x"01",x"20",x"0C",x"EE"
		,x"A9",x"01",x"A0",x"00",x"91",x"02",x"20",x"69"
		,x"DF",x"C9",x"00",x"F0",x"06",x"A2",x"00",x"8A"
		,x"4C",x"66",x"D4",x"A0",x"03",x"20",x"E9",x"EC"
		,x"A0",x"0B",x"20",x"49",x"E9",x"A0",x"1C",x"20"
		,x"E4",x"ED",x"A2",x"00",x"A9",x"01",x"A0",x"0A"
		,x"4C",x"37",x"E7",x"20",x"14",x"E8",x"AD",x"40"
		,x"A4",x"AE",x"41",x"A4",x"20",x"D1",x"EC",x"A0"
		,x"0D",x"20",x"49",x"E9",x"C9",x"02",x"8A",x"E9"
		,x"00",x"A5",x"04",x"E9",x"00",x"A5",x"05",x"E9"
		,x"00",x"B0",x"03",x"4C",x"8A",x"D6",x"A0",x"0D"
		,x"20",x"49",x"E9",x"20",x"28",x"EA",x"A0",x"05"
		,x"20",x"29",x"E9",x"A0",x"0F",x"20",x"32",x"E9"
		,x"20",x"5F",x"EC",x"D0",x"03",x"4C",x"8A",x"D6"
		,x"A0",x"01",x"20",x"29",x"E9",x"A0",x"13",x"20"
		,x"32",x"E9",x"A0",x"02",x"20",x"0C",x"EE",x"A0"
		,x"01",x"20",x"29",x"E9",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"B1",x"0A",x"C9",x"01",x"F0",x"11"
		,x"C9",x"02",x"D0",x"03",x"4C",x"EB",x"D5",x"C9"
		,x"03",x"D0",x"03",x"4C",x"3C",x"D6",x"4C",x"8A"
		,x"D6",x"A0",x"0B",x"20",x"29",x"E9",x"20",x"96"
		,x"EC",x"20",x"3D",x"ED",x"A0",x"06",x"20",x"DB"
		,x"ED",x"A0",x"05",x"20",x"49",x"E9",x"20",x"28"
		,x"EA",x"A0",x"0B",x"20",x"29",x"E9",x"8A",x"A2"
		,x"00",x"4A",x"A0",x"00",x"86",x"04",x"86",x"05"
		,x"20",x"91",x"E8",x"20",x"28",x"EA",x"20",x"EC"
		,x"D3",x"AA",x"D0",x"03",x"4C",x"8A",x"D6",x"A0"
		,x"01",x"20",x"29",x"E9",x"18",x"69",x"20",x"90"
		,x"01",x"E8",x"85",x"04",x"86",x"05",x"A0",x"07"
		,x"20",x"29",x"E9",x"A8",x"8A",x"29",x"01",x"AA"
		,x"98",x"18",x"65",x"04",x"85",x"04",x"8A",x"65"
		,x"05",x"AA",x"A5",x"04",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"A2",x"00",x"B1",x"0A",x"A0",x"08"
		,x"20",x"DB",x"ED",x"A0",x"07",x"20",x"29",x"E9"
		,x"18",x"69",x"01",x"90",x"01",x"E8",x"A0",x"06"
		,x"20",x"DB",x"ED",x"A0",x"05",x"20",x"49",x"E9"
		,x"20",x"28",x"EA",x"A0",x"0B",x"20",x"29",x"E9"
		,x"8A",x"A2",x"00",x"4A",x"A0",x"00",x"86",x"04"
		,x"86",x"05",x"20",x"91",x"E8",x"20",x"28",x"EA"
		,x"20",x"EC",x"D3",x"AA",x"D0",x"03",x"4C",x"8A"
		,x"D6",x"A0",x"09",x"20",x"29",x"E9",x"85",x"04"
		,x"86",x"05",x"A0",x"01",x"20",x"29",x"E9",x"18"
		,x"69",x"20",x"90",x"01",x"E8",x"85",x"0A",x"86"
		,x"0B",x"A0",x"07",x"20",x"29",x"E9",x"A8",x"8A"
		,x"29",x"01",x"AA",x"98",x"18",x"65",x"0A",x"85"
		,x"0A",x"8A",x"65",x"0B",x"AA",x"A5",x"0A",x"A0"
		,x"00",x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"AA"
		,x"98",x"05",x"04",x"85",x"04",x"8A",x"05",x"05"
		,x"AA",x"A5",x"04",x"A0",x"08",x"20",x"DB",x"ED"
		,x"A0",x"0D",x"20",x"49",x"E9",x"A2",x"00",x"86"
		,x"05",x"86",x"04",x"29",x"01",x"20",x"D0",x"EB"
		,x"F0",x"0B",x"A0",x"09",x"20",x"29",x"E9",x"20"
		,x"45",x"ED",x"4C",x"92",x"D6",x"A0",x"09",x"20"
		,x"29",x"E9",x"A8",x"8A",x"29",x"0F",x"AA",x"98"
		,x"4C",x"92",x"D6",x"A0",x"05",x"20",x"49",x"E9"
		,x"20",x"28",x"EA",x"A0",x"11",x"20",x"49",x"E9"
		,x"8A",x"A6",x"04",x"A4",x"05",x"84",x"04",x"A0"
		,x"00",x"84",x"05",x"20",x"91",x"E8",x"20",x"28"
		,x"EA",x"20",x"EC",x"D3",x"AA",x"F0",x"7B",x"A0"
		,x"01",x"20",x"29",x"E9",x"18",x"69",x"20",x"90"
		,x"01",x"E8",x"20",x"D1",x"EC",x"A0",x"0D",x"20"
		,x"29",x"E9",x"20",x"54",x"E7",x"A8",x"8A",x"29"
		,x"01",x"AA",x"98",x"20",x"1E",x"E7",x"A0",x"01"
		,x"20",x"1C",x"E9",x"A0",x"00",x"84",x"04",x"84"
		,x"05",x"4C",x"92",x"D6",x"A0",x"05",x"20",x"49"
		,x"E9",x"20",x"28",x"EA",x"A0",x"11",x"20",x"49"
		,x"E9",x"20",x"28",x"EA",x"A2",x"00",x"86",x"04"
		,x"86",x"05",x"A9",x"07",x"20",x"17",x"EB",x"20"
		,x"91",x"E8",x"20",x"28",x"EA",x"20",x"EC",x"D3"
		,x"AA",x"F0",x"27",x"A0",x"01",x"20",x"29",x"E9"
		,x"18",x"69",x"20",x"90",x"01",x"E8",x"20",x"D1"
		,x"EC",x"A0",x"0D",x"20",x"29",x"E9",x"20",x"5C"
		,x"E7",x"A8",x"8A",x"29",x"01",x"AA",x"98",x"20"
		,x"1E",x"E7",x"A0",x"03",x"20",x"32",x"E9",x"4C"
		,x"92",x"D6",x"A2",x"00",x"86",x"04",x"86",x"05"
		,x"A9",x"01",x"A0",x"0E",x"4C",x"37",x"E7",x"AD"
		,x"40",x"A4",x"AE",x"41",x"A4",x"20",x"D1",x"EC"
		,x"A2",x"00",x"86",x"04",x"86",x"05",x"A9",x"02"
		,x"A8",x"20",x"8A",x"EB",x"A0",x"05",x"20",x"49"
		,x"E9",x"20",x"28",x"EA",x"A0",x"05",x"20",x"29"
		,x"E9",x"A0",x"0F",x"20",x"32",x"E9",x"20",x"53"
		,x"EC",x"F0",x"0A",x"A2",x"00",x"86",x"04",x"86"
		,x"05",x"8A",x"4C",x"87",x"E8",x"A0",x"05",x"20"
		,x"49",x"E9",x"20",x"28",x"EA",x"A0",x"05",x"20"
		,x"29",x"E9",x"A0",x"02",x"85",x"0A",x"86",x"0B"
		,x"A2",x"00",x"B1",x"0A",x"86",x"04",x"86",x"05"
		,x"20",x"A8",x"E9",x"20",x"28",x"EA",x"A0",x"05"
		,x"20",x"29",x"E9",x"A0",x"1B",x"20",x"32",x"E9"
		,x"20",x"91",x"E8",x"4C",x"87",x"E8",x"AD",x"40"
		,x"A4",x"AE",x"41",x"A4",x"20",x"D1",x"EC",x"A0"
		,x"01",x"20",x"29",x"E9",x"18",x"69",x"20",x"90"
		,x"01",x"E8",x"20",x"D1",x"EC",x"A2",x"02",x"A9"
		,x"00",x"20",x"B9",x"E6",x"20",x"07",x"E8",x"A0"
		,x"08",x"20",x"29",x"E9",x"18",x"69",x"20",x"90"
		,x"01",x"E8",x"A0",x"05",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"A0",x"0C",x"20",x"49",x"E9",x"A0"
		,x"01",x"20",x"0C",x"EE",x"A9",x"01",x"A0",x"00"
		,x"91",x"02",x"20",x"69",x"DF",x"C9",x"00",x"F0"
		,x"03",x"4C",x"1A",x"D8",x"A0",x"01",x"20",x"29"
		,x"E9",x"18",x"69",x"1E",x"90",x"01",x"E8",x"E8"
		,x"E8",x"A0",x"01",x"20",x"1C",x"E9",x"E0",x"AA"
		,x"F0",x"03",x"4C",x"1A",x"D8",x"C9",x"55",x"F0"
		,x"03",x"4C",x"1A",x"D8",x"20",x"E0",x"E7",x"A0"
		,x"05",x"20",x"29",x"E9",x"18",x"69",x"56",x"90"
		,x"01",x"E8",x"A0",x"02",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"A9",x"A2",x"A2",x"EF",x"A0",x"00"
		,x"91",x"02",x"C8",x"8A",x"91",x"02",x"A2",x"00"
		,x"A9",x"05",x"20",x"43",x"E6",x"86",x"12",x"05"
		,x"12",x"D0",x"06",x"AA",x"A9",x"01",x"4C",x"87"
		,x"E8",x"20",x"E0",x"E7",x"A0",x"05",x"20",x"29"
		,x"E9",x"18",x"69",x"56",x"90",x"01",x"E8",x"A0"
		,x"02",x"91",x"02",x"C8",x"8A",x"91",x"02",x"A9"
		,x"A7",x"A2",x"EF",x"A0",x"00",x"91",x"02",x"C8"
		,x"8A",x"91",x"02",x"A2",x"00",x"A9",x"05",x"20"
		,x"43",x"E6",x"86",x"12",x"05",x"12",x"D0",x"06"
		,x"AA",x"A9",x"02",x"4C",x"87",x"E8",x"20",x"E0"
		,x"E7",x"A0",x"05",x"20",x"29",x"E9",x"18",x"69"
		,x"72",x"90",x"01",x"E8",x"A0",x"02",x"91",x"02"
		,x"C8",x"8A",x"91",x"02",x"A9",x"AC",x"A2",x"EF"
		,x"A0",x"00",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A2",x"00",x"A9",x"05",x"20",x"43",x"E6",x"86"
		,x"12",x"05",x"12",x"D0",x"15",x"A0",x"01",x"20"
		,x"29",x"E9",x"A0",x"48",x"85",x"0A",x"86",x"0B"
		,x"B1",x"0A",x"D0",x"06",x"AA",x"A9",x"03",x"4C"
		,x"87",x"E8",x"A2",x"00",x"8A",x"4C",x"87",x"E8"
		,x"20",x"FA",x"E7",x"AD",x"40",x"A4",x"AE",x"41"
		,x"A4",x"20",x"D1",x"EC",x"A0",x"09",x"20",x"29"
		,x"E9",x"A0",x"0D",x"20",x"1C",x"E9",x"18",x"69"
		,x"01",x"90",x"01",x"E8",x"A0",x"02",x"20",x"DB"
		,x"ED",x"29",x"0F",x"F0",x"03",x"4C",x"2E",x"D9"
		,x"A0",x"09",x"20",x"29",x"E9",x"20",x"D1",x"EC"
		,x"A0",x"0B",x"20",x"32",x"E9",x"20",x"40",x"EA"
		,x"A0",x"01",x"20",x"97",x"E9",x"A0",x"08",x"20"
		,x"E4",x"ED",x"20",x"4F",x"EA",x"A0",x"09",x"20"
		,x"29",x"E9",x"A0",x"07",x"20",x"32",x"E9",x"20"
		,x"CE",x"E8",x"F0",x"1D",x"A0",x"05",x"20",x"E9"
		,x"EC",x"A0",x"03",x"20",x"29",x"E9",x"A0",x"05"
		,x"20",x"1C",x"E9",x"20",x"2F",x"E8",x"B0",x"03"
		,x"4C",x"2E",x"D9",x"A2",x"00",x"8A",x"4C",x"48"
		,x"D9",x"A0",x"03",x"20",x"29",x"E9",x"20",x"45"
		,x"ED",x"85",x"0C",x"86",x"0D",x"A0",x"01",x"20"
		,x"29",x"E9",x"A0",x"02",x"85",x"0A",x"86",x"0B"
		,x"A2",x"00",x"B1",x"0A",x"38",x"E9",x"01",x"B0"
		,x"01",x"CA",x"25",x"0C",x"85",x"0C",x"8A",x"25"
		,x"0D",x"AA",x"A5",x"0C",x"E0",x"00",x"D0",x"6E"
		,x"C9",x"00",x"D0",x"6A",x"A0",x"09",x"20",x"29"
		,x"E9",x"A0",x"07",x"20",x"32",x"E9",x"20",x"28"
		,x"EA",x"20",x"6B",x"D4",x"A0",x"04",x"20",x"0C"
		,x"EE",x"A0",x"07",x"20",x"49",x"E9",x"20",x"28"
		,x"EA",x"A0",x"05",x"20",x"29",x"E9",x"A0",x"0F"
		,x"20",x"32",x"E9",x"20",x"53",x"EC",x"D0",x"14"
		,x"A0",x"07",x"20",x"49",x"E9",x"C9",x"02",x"8A"
		,x"E9",x"00",x"A5",x"04",x"E9",x"00",x"A5",x"05"
		,x"E9",x"00",x"B0",x"06",x"A2",x"00",x"8A",x"4C"
		,x"48",x"D9",x"A0",x"0B",x"20",x"E9",x"EC",x"A0"
		,x"09",x"20",x"49",x"E9",x"A0",x"04",x"20",x"E4"
		,x"ED",x"A0",x"0B",x"20",x"E9",x"EC",x"A0",x"09"
		,x"20",x"49",x"E9",x"20",x"28",x"EA",x"20",x"97"
		,x"D6",x"A0",x"08",x"20",x"E4",x"ED",x"A0",x"09"
		,x"20",x"29",x"E9",x"85",x"04",x"86",x"05",x"A0"
		,x"03",x"20",x"29",x"E9",x"A0",x"0C",x"91",x"04"
		,x"C8",x"8A",x"91",x"04",x"A2",x"00",x"A9",x"01"
		,x"A0",x"0A",x"4C",x"37",x"E7",x"20",x"ED",x"E7"
		,x"A0",x"08",x"20",x"E9",x"EC",x"A2",x"00",x"A9"
		,x"20",x"20",x"D1",x"EC",x"A9",x"0B",x"20",x"C1"
		,x"E6",x"A9",x"00",x"A0",x"01",x"91",x"02",x"A9"
		,x"18",x"88",x"91",x"02",x"98",x"A0",x"04",x"91"
		,x"02",x"A9",x"08",x"88",x"91",x"02",x"A0",x"08"
		,x"20",x"29",x"E9",x"85",x"0C",x"86",x"0D",x"A0"
		,x"01",x"20",x"1C",x"E9",x"85",x"06",x"86",x"07"
		,x"18",x"69",x"01",x"90",x"01",x"E8",x"A0",x"00"
		,x"91",x"0C",x"C8",x"8A",x"91",x"0C",x"88",x"B1"
		,x"06",x"A0",x"02",x"91",x"02",x"C9",x"21",x"B0"
		,x"04",x"A9",x"00",x"91",x"02",x"B1",x"02",x"F0"
		,x"06",x"B1",x"02",x"C9",x"2F",x"D0",x"26",x"A0"
		,x"04",x"B1",x"02",x"D0",x"03",x"4C",x"1F",x"DB"
		,x"A0",x"06",x"20",x"29",x"E9",x"85",x"04",x"86"
		,x"05",x"A2",x"00",x"A0",x"00",x"B1",x"02",x"C8"
		,x"31",x"02",x"A0",x"0B",x"91",x"04",x"A0",x"02"
		,x"B1",x"02",x"4C",x"23",x"DB",x"B1",x"02",x"C9"
		,x"2E",x"D0",x"27",x"88",x"B1",x"02",x"29",x"01"
		,x"F0",x"03",x"4C",x"1F",x"DB",x"A0",x"04",x"B1"
		,x"02",x"C9",x"01",x"B0",x"03",x"4C",x"1F",x"DB"
		,x"B1",x"02",x"C9",x"09",x"90",x"03",x"4C",x"1F"
		,x"DB",x"A9",x"08",x"91",x"02",x"A9",x"0B",x"4C"
		,x"73",x"D9",x"B1",x"02",x"C9",x"81",x"90",x"06"
		,x"B1",x"02",x"C9",x"A0",x"90",x"0C",x"B1",x"02"
		,x"C9",x"E0",x"90",x"21",x"B1",x"02",x"C9",x"FD"
		,x"B0",x"1B",x"A0",x"04",x"B1",x"02",x"D0",x"0C"
		,x"A0",x"02",x"B1",x"02",x"C9",x"E5",x"D0",x"04"
		,x"A9",x"05",x"91",x"02",x"A0",x"01",x"B1",x"02"
		,x"49",x"01",x"4C",x"E5",x"DA",x"B1",x"02",x"C9"
		,x"7F",x"90",x"09",x"B1",x"02",x"C9",x"81",x"B0"
		,x"03",x"4C",x"1F",x"DB",x"B1",x"02",x"C9",x"22"
		,x"D0",x"03",x"4C",x"1F",x"DB",x"B1",x"02",x"C9"
		,x"2A",x"B0",x"03",x"4C",x"DF",x"DA",x"B1",x"02"
		,x"C9",x"2D",x"B0",x"03",x"4C",x"1F",x"DB",x"B1"
		,x"02",x"C9",x"3A",x"90",x"7A",x"B1",x"02",x"C9"
		,x"40",x"B0",x"03",x"4C",x"1F",x"DB",x"88",x"B1"
		,x"02",x"29",x"01",x"D0",x"6A",x"C8",x"B1",x"02"
		,x"C9",x"7C",x"D0",x"03",x"4C",x"1F",x"DB",x"B1"
		,x"02",x"C9",x"5B",x"90",x"09",x"B1",x"02",x"C9"
		,x"5E",x"B0",x"03",x"4C",x"1F",x"DB",x"B1",x"02"
		,x"C9",x"41",x"90",x"1E",x"B1",x"02",x"C9",x"5B"
		,x"B0",x"18",x"C8",x"B1",x"02",x"C9",x"08",x"D0"
		,x"09",x"A0",x"00",x"B1",x"02",x"29",x"F7",x"4C"
		,x"B0",x"DA",x"A0",x"00",x"B1",x"02",x"29",x"EF"
		,x"91",x"02",x"A0",x"02",x"B1",x"02",x"C9",x"61"
		,x"90",x"25",x"B1",x"02",x"C9",x"7B",x"B0",x"1F"
		,x"38",x"B1",x"02",x"E9",x"20",x"91",x"02",x"C8"
		,x"B1",x"02",x"C9",x"08",x"D0",x"09",x"A0",x"01"
		,x"B1",x"02",x"09",x"08",x"4C",x"DD",x"DA",x"A0"
		,x"01",x"B1",x"02",x"09",x"10",x"91",x"02",x"A0"
		,x"01",x"B1",x"02",x"29",x"FE",x"91",x"02",x"A0"
		,x"04",x"A2",x"00",x"B1",x"02",x"20",x"D1",x"EC"
		,x"A0",x"05",x"B1",x"02",x"20",x"2F",x"E8",x"B0"
		,x"26",x"A0",x"04",x"B1",x"02",x"48",x"18",x"69"
		,x"01",x"91",x"02",x"68",x"C8",x"18",x"71",x"02"
		,x"48",x"A9",x"00",x"C8",x"71",x"02",x"AA",x"68"
		,x"85",x"0A",x"86",x"0B",x"A0",x"02",x"B1",x"02"
		,x"A0",x"00",x"91",x"0A",x"4C",x"76",x"D9",x"A2"
		,x"00",x"A9",x"01",x"A0",x"09",x"4C",x"37",x"E7"
		,x"20",x"ED",x"E7",x"A2",x"00",x"8A",x"20",x"D1"
		,x"EC",x"AD",x"40",x"A4",x"AE",x"41",x"A4",x"20"
		,x"D1",x"EC",x"A0",x"01",x"20",x"29",x"E9",x"A0"
		,x"17",x"20",x"32",x"E9",x"A0",x"05",x"20",x"0C"
		,x"EE",x"A0",x"01",x"20",x"29",x"E9",x"A0",x"00"
		,x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"C9",x"03"
		,x"D0",x"2C",x"A0",x"12",x"20",x"E9",x"EC",x"A0"
		,x"14",x"20",x"E9",x"EC",x"A0",x"0C",x"20",x"49"
		,x"E9",x"A0",x"00",x"20",x"E4",x"ED",x"A0",x"04"
		,x"20",x"E4",x"ED",x"A0",x"12",x"20",x"E9",x"EC"
		,x"A0",x"0A",x"20",x"49",x"E9",x"20",x"28",x"EA"
		,x"20",x"97",x"D6",x"4C",x"AA",x"DB",x"A0",x"12"
		,x"20",x"E9",x"EC",x"A0",x"14",x"20",x"E9",x"EC"
		,x"A2",x"00",x"86",x"04",x"86",x"05",x"8A",x"A8"
		,x"20",x"E4",x"ED",x"A0",x"04",x"20",x"E4",x"ED"
		,x"A0",x"12",x"20",x"E9",x"EC",x"A0",x"0A",x"20"
		,x"49",x"E9",x"A0",x"08",x"20",x"E4",x"ED",x"A0"
		,x"10",x"20",x"29",x"E9",x"85",x"0A",x"86",x"0B"
		,x"A9",x"00",x"A0",x"0C",x"91",x"0A",x"C8",x"91"
		,x"0A",x"A0",x"0C",x"20",x"29",x"E9",x"A0",x"00"
		,x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"C9",x"20"
		,x"F0",x"11",x"A0",x"0C",x"20",x"29",x"E9",x"A0"
		,x"00",x"85",x"0A",x"86",x"0B",x"B1",x"0A",x"C9"
		,x"2F",x"D0",x"13",x"A0",x"0C",x"20",x"29",x"E9"
		,x"18",x"69",x"01",x"90",x"01",x"E8",x"A0",x"0B"
		,x"20",x"DB",x"ED",x"4C",x"C1",x"DB",x"A0",x"0C"
		,x"20",x"29",x"E9",x"A0",x"00",x"85",x"0A",x"86"
		,x"0B",x"B1",x"0A",x"C9",x"20",x"B0",x"15",x"A0"
		,x"0A",x"20",x"29",x"E9",x"85",x"04",x"86",x"05"
		,x"A9",x"00",x"A8",x"91",x"04",x"C8",x"91",x"04"
		,x"AA",x"4C",x"D9",x"DD",x"20",x"E0",x"E7",x"A9"
		,x"0F",x"18",x"A6",x"03",x"65",x"02",x"90",x"01"
		,x"E8",x"A0",x"02",x"91",x"02",x"C8",x"8A",x"91"
		,x"02",x"A0",x"12",x"20",x"29",x"E9",x"A0",x"00"
		,x"91",x"02",x"C8",x"8A",x"91",x"02",x"20",x"4D"
		,x"D9",x"A0",x"04",x"91",x"02",x"C9",x"01",x"D0"
		,x"06",x"A2",x"00",x"98",x"4C",x"D9",x"DD",x"A0"
		,x"10",x"20",x"29",x"E9",x"A0",x"0B",x"20",x"32"
		,x"E9",x"20",x"28",x"EA",x"20",x"EC",x"D3",x"AA"
		,x"D0",x"05",x"A9",x"07",x"4C",x"D9",x"DD",x"A0"
		,x"01",x"20",x"29",x"E9",x"18",x"69",x"20",x"90"
		,x"01",x"E8",x"20",x"D1",x"EC",x"A0",x"12",x"20"
		,x"29",x"E9",x"A0",x"0D",x"20",x"1C",x"E9",x"A2"
		,x"00",x"29",x"0F",x"20",x"D1",x"EC",x"A9",x"05"
		,x"20",x"07",x"ED",x"20",x"1E",x"E7",x"A0",x"02"
		,x"20",x"DB",x"ED",x"A0",x"00",x"85",x"0A",x"86"
		,x"0B",x"B1",x"0A",x"D0",x"13",x"A0",x"04",x"B1"
		,x"02",x"D0",x"06",x"AA",x"A9",x"02",x"4C",x"D9"
		,x"DD",x"A2",x"00",x"A9",x"03",x"4C",x"D9",x"DD"
		,x"A0",x"03",x"20",x"29",x"E9",x"A0",x"00",x"85"
		,x"0A",x"86",x"0B",x"B1",x"0A",x"C9",x"E5",x"F0"
		,x"41",x"A0",x"03",x"20",x"29",x"E9",x"18",x"69"
		,x"0B",x"90",x"01",x"E8",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"B1",x"0A",x"29",x"08",x"D0",x"2A"
		,x"20",x"E0",x"E7",x"A0",x"07",x"20",x"29",x"E9"
		,x"A0",x"02",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A0",x"12",x"20",x"29",x"E9",x"A0",x"00",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"A2",x"00",x"A9"
		,x"0B",x"20",x"43",x"E6",x"86",x"12",x"05",x"12"
		,x"F0",x"1E",x"A0",x"12",x"20",x"E9",x"EC",x"20"
		,x"20",x"D8",x"AA",x"F0",x"03",x"4C",x"4F",x"DC"
		,x"A0",x"04",x"B1",x"02",x"D0",x"05",x"A9",x"02"
		,x"4C",x"D9",x"DD",x"A9",x"03",x"4C",x"D9",x"DD"
		,x"A0",x"04",x"B1",x"02",x"D0",x"1C",x"A0",x"0A"
		,x"20",x"29",x"E9",x"85",x"04",x"86",x"05",x"A0"
		,x"03",x"20",x"29",x"E9",x"A0",x"00",x"91",x"04"
		,x"C8",x"8A",x"91",x"04",x"A2",x"00",x"8A",x"4C"
		,x"D9",x"DD",x"88",x"20",x"29",x"E9",x"18",x"69"
		,x"0B",x"90",x"01",x"E8",x"A0",x"00",x"85",x"0A"
		,x"86",x"0B",x"B1",x"0A",x"29",x"10",x"D0",x"06"
		,x"AA",x"A9",x"03",x"4C",x"D9",x"DD",x"A0",x"03"
		,x"20",x"29",x"E9",x"18",x"69",x"14",x"90",x"01"
		,x"E8",x"A0",x"01",x"20",x"1C",x"E9",x"86",x"05"
		,x"85",x"04",x"A9",x"00",x"AA",x"20",x"28",x"EA"
		,x"A0",x"07",x"20",x"29",x"E9",x"18",x"69",x"1A"
		,x"90",x"01",x"E8",x"A0",x"01",x"20",x"1C",x"E9"
		,x"A0",x"00",x"84",x"04",x"84",x"05",x"20",x"04"
		,x"EA",x"A0",x"05",x"20",x"0C",x"EE",x"A0",x"12"
		,x"20",x"E9",x"EC",x"A0",x"14",x"20",x"E9",x"EC"
		,x"A0",x"0C",x"20",x"49",x"E9",x"A0",x"00",x"20"
		,x"E4",x"ED",x"A0",x"04",x"20",x"E4",x"ED",x"A0"
		,x"12",x"20",x"E9",x"EC",x"A0",x"0A",x"20",x"49"
		,x"E9",x"20",x"28",x"EA",x"20",x"97",x"D6",x"A0"
		,x"08",x"20",x"E4",x"ED",x"A0",x"10",x"20",x"29"
		,x"E9",x"85",x"04",x"86",x"05",x"A9",x"00",x"A0"
		,x"0C",x"91",x"04",x"C8",x"91",x"04",x"4C",x"1C"
		,x"DC",x"A0",x"11",x"4C",x"37",x"E7",x"20",x"21"
		,x"E8",x"AD",x"40",x"A4",x"AE",x"41",x"A4",x"20"
		,x"D1",x"EC",x"A0",x"01",x"B1",x"02",x"88",x"11"
		,x"02",x"D0",x"06",x"AA",x"A9",x"0A",x"4C",x"35"
		,x"DE",x"20",x"63",x"DF",x"29",x"01",x"F0",x"1C"
		,x"A0",x"01",x"20",x"29",x"E9",x"A0",x"01",x"85"
		,x"0A",x"86",x"0B",x"B1",x"0A",x"F0",x"07",x"A2"
		,x"00",x"A9",x"08",x"4C",x"35",x"DE",x"20",x"6C"
		,x"D1",x"4C",x"35",x"DE",x"A0",x"01",x"20",x"29"
		,x"E9",x"A0",x"00",x"85",x"0A",x"86",x"0B",x"B1"
		,x"0A",x"AA",x"D0",x"06",x"20",x"6C",x"D1",x"4C"
		,x"35",x"DE",x"A2",x"00",x"8A",x"A0",x"02",x"4C"
		,x"7E",x"E9",x"20",x"C6",x"E7",x"A9",x"01",x"8D"
		,x"02",x"B5",x"A9",x"00",x"8D",x"00",x"A0",x"A8"
		,x"91",x"02",x"AD",x"00",x"A0",x"29",x"02",x"F0"
		,x"03",x"4C",x"37",x"DF",x"A9",x"0A",x"C8",x"91"
		,x"02",x"20",x"91",x"E3",x"A0",x"01",x"38",x"B1"
		,x"02",x"E9",x"01",x"91",x"02",x"AA",x"D0",x"F1"
		,x"8D",x"02",x"B5",x"20",x"ED",x"E7",x"A9",x"40"
		,x"A0",x"04",x"91",x"02",x"A0",x"00",x"8A",x"91"
		,x"02",x"C8",x"91",x"02",x"C8",x"91",x"02",x"C8"
		,x"91",x"02",x"20",x"0A",x"E5",x"C9",x"01",x"D0"
		,x"78",x"A9",x"32",x"8D",x"42",x"A4",x"AD",x"42"
		,x"A4",x"F0",x"1D",x"20",x"ED",x"E7",x"A9",x"41"
		,x"A0",x"04",x"91",x"02",x"A0",x"00",x"98",x"91"
		,x"02",x"C8",x"91",x"02",x"C8",x"91",x"02",x"C8"
		,x"91",x"02",x"20",x"0A",x"E5",x"AA",x"D0",x"DE"
		,x"AD",x"42",x"A4",x"D0",x"46",x"A9",x"64",x"8D"
		,x"42",x"A4",x"AD",x"42",x"A4",x"F0",x"42",x"20"
		,x"ED",x"E7",x"A9",x"77",x"A0",x"04",x"91",x"02"
		,x"A0",x"00",x"98",x"91",x"02",x"C8",x"91",x"02"
		,x"C8",x"91",x"02",x"C8",x"91",x"02",x"20",x"0A"
		,x"E5",x"29",x"FE",x"D0",x"DD",x"20",x"ED",x"E7"
		,x"A9",x"69",x"A0",x"04",x"91",x"02",x"A0",x"00"
		,x"98",x"91",x"02",x"C8",x"91",x"02",x"C8",x"91"
		,x"02",x"C8",x"91",x"02",x"20",x"0A",x"E5",x"C9"
		,x"00",x"D0",x"BF",x"A9",x"01",x"A0",x"00",x"91"
		,x"02",x"A0",x"00",x"B1",x"02",x"F0",x"28",x"20"
		,x"ED",x"E7",x"A9",x"50",x"A0",x"04",x"91",x"02"
		,x"A9",x"00",x"A8",x"91",x"02",x"A0",x"02",x"91"
		,x"02",x"C8",x"91",x"02",x"A9",x"02",x"A0",x"01"
		,x"91",x"02",x"20",x"0A",x"E5",x"C9",x"00",x"D0"
		,x"06",x"A9",x"02",x"A0",x"00",x"91",x"02",x"A9"
		,x"01",x"8D",x"02",x"B5",x"20",x"91",x"E3",x"A0"
		,x"00",x"B1",x"02",x"C9",x"02",x"D0",x"0B",x"AD"
		,x"00",x"A0",x"29",x"FE",x"8D",x"00",x"A0",x"4C"
		,x"4D",x"DF",x"20",x"55",x"DF",x"A2",x"00",x"AD"
		,x"00",x"A0",x"4C",x"6A",x"E8",x"AD",x"00",x"A0"
		,x"09",x"01",x"8D",x"00",x"A0",x"A2",x"00",x"AD"
		,x"00",x"A0",x"60",x"A2",x"00",x"AD",x"00",x"A0"
		,x"60",x"AD",x"00",x"A0",x"29",x"01",x"F0",x"07"
		,x"A2",x"00",x"A9",x"03",x"4C",x"8C",x"E8",x"A8"
		,x"B1",x"02",x"D0",x"06",x"AA",x"A9",x"04",x"4C"
		,x"8C",x"E8",x"A0",x"04",x"20",x"49",x"E9",x"20"
		,x"28",x"EA",x"A2",x"00",x"86",x"04",x"86",x"05"
		,x"A9",x"09",x"20",x"5C",x"EA",x"A0",x"01",x"20"
		,x"0C",x"EE",x"A9",x"00",x"8D",x"02",x"B5",x"A8"
		,x"B1",x"02",x"C9",x"01",x"D0",x"40",x"20",x"ED"
		,x"E7",x"A9",x"51",x"A0",x"04",x"91",x"02",x"A0"
		,x"09",x"20",x"49",x"E9",x"A0",x"00",x"20",x"0C"
		,x"EE",x"20",x"0A",x"E5",x"C9",x"00",x"F0",x"03"
		,x"4C",x"51",x"E0",x"20",x"D3",x"E7",x"A0",x"09"
		,x"20",x"29",x"E9",x"A0",x"01",x"91",x"02",x"C8"
		,x"8A",x"91",x"02",x"A9",x"00",x"A8",x"91",x"02"
		,x"20",x"C4",x"E3",x"AA",x"F0",x"73",x"A9",x"00"
		,x"A8",x"91",x"02",x"4C",x"51",x"E0",x"20",x"ED"
		,x"E7",x"A9",x"52",x"A0",x"04",x"91",x"02",x"A0"
		,x"09",x"20",x"49",x"E9",x"A0",x"00",x"20",x"0C"
		,x"EE",x"20",x"0A",x"E5",x"C9",x"00",x"D0",x"51"
		,x"20",x"D3",x"E7",x"A0",x"09",x"20",x"29",x"E9"
		,x"A0",x"01",x"91",x"02",x"C8",x"8A",x"91",x"02"
		,x"A9",x"00",x"A8",x"91",x"02",x"20",x"C4",x"E3"
		,x"AA",x"F0",x"1C",x"A0",x"05",x"18",x"A9",x"00"
		,x"71",x"02",x"91",x"02",x"C8",x"A9",x"02",x"71"
		,x"02",x"91",x"02",x"A0",x"00",x"38",x"B1",x"02"
		,x"E9",x"01",x"91",x"02",x"AA",x"D0",x"C9",x"20"
		,x"ED",x"E7",x"A9",x"4C",x"A0",x"04",x"91",x"02"
		,x"A0",x"00",x"8A",x"91",x"02",x"C8",x"91",x"02"
		,x"C8",x"91",x"02",x"C8",x"91",x"02",x"20",x"0A"
		,x"E5",x"A9",x"01",x"8D",x"02",x"B5",x"20",x"91"
		,x"E3",x"A0",x"00",x"B1",x"02",x"F0",x"07",x"A2"
		,x"00",x"A9",x"01",x"4C",x"8C",x"E8",x"AA",x"4C"
		,x"8C",x"E8",x"AD",x"00",x"A0",x"29",x"01",x"F0"
		,x"07",x"A2",x"00",x"A9",x"03",x"4C",x"8C",x"E8"
		,x"AD",x"00",x"A0",x"29",x"04",x"F0",x"07",x"A2"
		,x"00",x"A9",x"02",x"4C",x"8C",x"E8",x"A8",x"B1"
		,x"02",x"D0",x"06",x"AA",x"A9",x"04",x"4C",x"8C"
		,x"E8",x"A0",x"04",x"20",x"49",x"E9",x"20",x"28"
		,x"EA",x"A2",x"00",x"86",x"04",x"86",x"05",x"A9"
		,x"09",x"20",x"5C",x"EA",x"A0",x"01",x"20",x"0C"
		,x"EE",x"A9",x"00",x"8D",x"02",x"B5",x"A8",x"B1"
		,x"02",x"C9",x"01",x"D0",x"3E",x"20",x"ED",x"E7"
		,x"A9",x"58",x"A0",x"04",x"91",x"02",x"A0",x"09"
		,x"20",x"49",x"E9",x"A0",x"00",x"20",x"0C",x"EE"
		,x"20",x"0A",x"E5",x"C9",x"00",x"F0",x"03",x"4C"
		,x"62",x"E1",x"20",x"D3",x"E7",x"A0",x"09",x"20"
		,x"29",x"E9",x"A0",x"01",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"A9",x"FE",x"A0",x"00",x"91",x"02"
		,x"20",x"5E",x"E4",x"AA",x"F0",x"74",x"A9",x"00"
		,x"4C",x"5E",x"E1",x"20",x"ED",x"E7",x"A9",x"59"
		,x"A0",x"04",x"91",x"02",x"A0",x"09",x"20",x"49"
		,x"E9",x"A0",x"00",x"20",x"0C",x"EE",x"20",x"0A"
		,x"E5",x"C9",x"00",x"D0",x"55",x"20",x"D3",x"E7"
		,x"A0",x"09",x"20",x"29",x"E9",x"A0",x"01",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"A9",x"FC",x"A0"
		,x"00",x"91",x"02",x"20",x"5E",x"E4",x"AA",x"F0"
		,x"1C",x"A0",x"05",x"18",x"A9",x"00",x"71",x"02"
		,x"91",x"02",x"C8",x"A9",x"02",x"71",x"02",x"91"
		,x"02",x"A0",x"00",x"38",x"B1",x"02",x"E9",x"01"
		,x"91",x"02",x"AA",x"D0",x"C8",x"20",x"D3",x"E7"
		,x"8A",x"A0",x"01",x"91",x"02",x"C8",x"91",x"02"
		,x"A9",x"FD",x"A0",x"00",x"91",x"02",x"20",x"5E"
		,x"E4",x"AA",x"D0",x"06",x"A9",x"01",x"A0",x"00"
		,x"91",x"02",x"A9",x"01",x"8D",x"02",x"B5",x"20"
		,x"91",x"E3",x"A0",x"00",x"B1",x"02",x"F0",x"07"
		,x"A2",x"00",x"A9",x"01",x"4C",x"8C",x"E8",x"AA"
		,x"4C",x"8C",x"E8",x"A0",x"12",x"20",x"49",x"EE"
		,x"A0",x"15",x"20",x"E9",x"EC",x"20",x"E0",x"E7"
		,x"AD",x"00",x"A0",x"29",x"01",x"F0",x"07",x"A2"
		,x"00",x"A9",x"03",x"4C",x"8C",x"E3",x"8D",x"02"
		,x"B5",x"A9",x"01",x"A0",x"17",x"91",x"02",x"A0"
		,x"1A",x"B1",x"02",x"C9",x"01",x"F0",x"18",x"C9"
		,x"0A",x"D0",x"03",x"4C",x"99",x"E2",x"C9",x"0B"
		,x"D0",x"03",x"4C",x"DE",x"E2",x"C9",x"0C",x"D0"
		,x"03",x"4C",x"20",x"E3",x"4C",x"78",x"E3",x"20"
		,x"ED",x"E7",x"A9",x"49",x"A0",x"04",x"91",x"02"
		,x"A0",x"00",x"98",x"91",x"02",x"C8",x"91",x"02"
		,x"C8",x"91",x"02",x"C8",x"91",x"02",x"20",x"0A"
		,x"E5",x"C9",x"00",x"F0",x"03",x"4C",x"7E",x"E3"
		,x"20",x"D3",x"E7",x"A9",x"09",x"18",x"A6",x"03"
		,x"65",x"02",x"90",x"01",x"E8",x"A0",x"01",x"91"
		,x"02",x"C8",x"8A",x"91",x"02",x"A9",x"08",x"A0"
		,x"00",x"91",x"02",x"20",x"C4",x"E3",x"AA",x"D0"
		,x"03",x"4C",x"7E",x"E3",x"A2",x"00",x"A9",x"01"
		,x"20",x"D1",x"EC",x"A0",x"12",x"B1",x"02",x"29"
		,x"80",x"20",x"D1",x"EC",x"A9",x"07",x"20",x"97"
		,x"ED",x"20",x"D1",x"EC",x"A0",x"13",x"B1",x"02"
		,x"A2",x"00",x"29",x"03",x"20",x"54",x"E7",x"20"
		,x"1E",x"E7",x"18",x"69",x"02",x"90",x"01",x"E8"
		,x"20",x"09",x"ED",x"A0",x"02",x"20",x"DB",x"ED"
		,x"A0",x"0E",x"B1",x"02",x"A2",x"00",x"29",x"03"
		,x"20",x"D1",x"EC",x"A9",x"06",x"20",x"97",x"ED"
		,x"20",x"D1",x"EC",x"A0",x"0F",x"A2",x"00",x"B1"
		,x"02",x"20",x"5C",x"E7",x"20",x"1E",x"E7",x"20"
		,x"D1",x"EC",x"A0",x"0E",x"B1",x"02",x"29",x"03"
		,x"AA",x"A9",x"00",x"20",x"5C",x"E7",x"20",x"1E"
		,x"E7",x"18",x"69",x"01",x"90",x"01",x"E8",x"A0"
		,x"00",x"20",x"DB",x"ED",x"A0",x"07",x"20",x"E9"
		,x"EC",x"A0",x"03",x"20",x"29",x"E9",x"A0",x"00"
		,x"84",x"04",x"84",x"05",x"20",x"28",x"EA",x"A0"
		,x"09",x"20",x"29",x"E9",x"20",x"A8",x"E9",x"A0"
		,x"00",x"20",x"E4",x"ED",x"A9",x"00",x"4C",x"7A"
		,x"E3",x"20",x"ED",x"E7",x"A9",x"49",x"A0",x"04"
		,x"91",x"02",x"A0",x"00",x"98",x"91",x"02",x"C8"
		,x"91",x"02",x"C8",x"91",x"02",x"C8",x"91",x"02"
		,x"20",x"0A",x"E5",x"C9",x"00",x"F0",x"03",x"4C"
		,x"7E",x"E3",x"20",x"D3",x"E7",x"A0",x"08",x"20"
		,x"29",x"E9",x"A0",x"01",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"A9",x"08",x"A0",x"00",x"91",x"02"
		,x"20",x"C4",x"E3",x"AA",x"D0",x"03",x"4C",x"7E"
		,x"E3",x"A9",x"00",x"4C",x"7A",x"E3",x"20",x"ED"
		,x"E7",x"A9",x"4A",x"A0",x"04",x"91",x"02",x"A0"
		,x"00",x"98",x"91",x"02",x"C8",x"91",x"02",x"C8"
		,x"91",x"02",x"C8",x"91",x"02",x"20",x"0A",x"E5"
		,x"C9",x"00",x"F0",x"03",x"4C",x"7E",x"E3",x"20"
		,x"D3",x"E7",x"A0",x"08",x"20",x"29",x"E9",x"A0"
		,x"01",x"91",x"02",x"C8",x"8A",x"91",x"02",x"A9"
		,x"08",x"A0",x"00",x"91",x"02",x"20",x"C4",x"E3"
		,x"AA",x"F0",x"63",x"A9",x"00",x"4C",x"7A",x"E3"
		,x"20",x"ED",x"E7",x"A9",x"7A",x"A0",x"04",x"91"
		,x"02",x"A0",x"00",x"98",x"91",x"02",x"C8",x"91"
		,x"02",x"C8",x"91",x"02",x"C8",x"91",x"02",x"20"
		,x"0A",x"E5",x"C9",x"00",x"D0",x"40",x"A0",x"16"
		,x"91",x"02",x"C9",x"04",x"B0",x"2D",x"A0",x"05"
		,x"20",x"29",x"E9",x"85",x"06",x"86",x"07",x"18"
		,x"69",x"01",x"90",x"01",x"E8",x"A0",x"04",x"20"
		,x"DB",x"ED",x"A5",x"06",x"A6",x"07",x"20",x"D1"
		,x"EC",x"20",x"91",x"E3",x"A0",x"00",x"20",x"C3"
		,x"ED",x"A0",x"16",x"B1",x"02",x"18",x"69",x"01"
		,x"4C",x"40",x"E3",x"A9",x"00",x"4C",x"7A",x"E3"
		,x"A9",x"04",x"A0",x"17",x"91",x"02",x"A9",x"01"
		,x"8D",x"02",x"B5",x"20",x"91",x"E3",x"A0",x"17"
		,x"A2",x"00",x"B1",x"02",x"A0",x"1B",x"4C",x"37"
		,x"E7",x"A9",x"FF",x"8D",x"00",x"B5",x"AD",x"01"
		,x"B5",x"29",x"01",x"D0",x"F9",x"AA",x"AD",x"00"
		,x"B5",x"60",x"20",x"BD",x"E7",x"A9",x"32",x"8D"
		,x"43",x"A4",x"20",x"91",x"E3",x"20",x"91",x"E3"
		,x"A0",x"00",x"91",x"02",x"C9",x"FF",x"F0",x"05"
		,x"AD",x"43",x"A4",x"D0",x"F0",x"A2",x"00",x"B1"
		,x"02",x"4C",x"5B",x"E8",x"20",x"BD",x"E7",x"A9"
		,x"0A",x"8D",x"42",x"A4",x"20",x"91",x"E3",x"A0"
		,x"00",x"91",x"02",x"C9",x"FF",x"D0",x"05",x"AD"
		,x"42",x"A4",x"D0",x"F0",x"B1",x"02",x"C9",x"FE"
		,x"F0",x"06",x"A2",x"00",x"8A",x"4C",x"7D",x"E8"
		,x"A9",x"FF",x"8D",x"00",x"B5",x"AD",x"01",x"B5"
		,x"29",x"01",x"D0",x"F9",x"A0",x"03",x"20",x"29"
		,x"E9",x"85",x"06",x"86",x"07",x"18",x"69",x"01"
		,x"90",x"01",x"E8",x"A0",x"02",x"20",x"DB",x"ED"
		,x"A5",x"06",x"A6",x"07",x"85",x"04",x"86",x"05"
		,x"AD",x"00",x"B5",x"A0",x"00",x"91",x"04",x"A9"
		,x"FF",x"8D",x"00",x"B5",x"AD",x"01",x"B5",x"29"
		,x"01",x"D0",x"F9",x"A0",x"03",x"20",x"29",x"E9"
		,x"85",x"06",x"86",x"07",x"18",x"69",x"01",x"90"
		,x"01",x"E8",x"A0",x"02",x"20",x"DB",x"ED",x"A5"
		,x"06",x"A6",x"07",x"85",x"04",x"86",x"05",x"AD"
		,x"00",x"B5",x"A0",x"00",x"91",x"04",x"C8",x"38"
		,x"B1",x"02",x"E9",x"01",x"91",x"02",x"AA",x"D0"
		,x"97",x"20",x"91",x"E3",x"20",x"91",x"E3",x"A2"
		,x"00",x"A9",x"01",x"4C",x"7D",x"E8",x"20",x"BD"
		,x"E7",x"A9",x"00",x"20",x"BB",x"EC",x"20",x"A2"
		,x"E3",x"C9",x"FF",x"F0",x"06",x"A2",x"00",x"8A"
		,x"4C",x"82",x"E8",x"A0",x"02",x"B1",x"02",x"8D"
		,x"00",x"B5",x"AD",x"01",x"B5",x"29",x"01",x"D0"
		,x"F9",x"A0",x"02",x"B1",x"02",x"C9",x"FD",x"F0"
		,x"7A",x"A0",x"04",x"20",x"29",x"E9",x"85",x"06"
		,x"86",x"07",x"18",x"69",x"01",x"90",x"01",x"E8"
		,x"A0",x"03",x"20",x"DB",x"ED",x"A0",x"00",x"B1"
		,x"06",x"8D",x"00",x"B5",x"AD",x"01",x"B5",x"29"
		,x"01",x"D0",x"F9",x"A0",x"04",x"20",x"29",x"E9"
		,x"85",x"06",x"86",x"07",x"18",x"69",x"01",x"90"
		,x"01",x"E8",x"A0",x"03",x"20",x"DB",x"ED",x"A0"
		,x"00",x"B1",x"06",x"8D",x"00",x"B5",x"AD",x"01"
		,x"B5",x"29",x"01",x"D0",x"F9",x"A8",x"38",x"B1"
		,x"02",x"E9",x"01",x"91",x"02",x"AA",x"D0",x"B1"
		,x"A9",x"FF",x"8D",x"00",x"B5",x"AD",x"01",x"B5"
		,x"29",x"01",x"D0",x"F9",x"A9",x"FF",x"8D",x"00"
		,x"B5",x"AD",x"01",x"B5",x"29",x"01",x"D0",x"F9"
		,x"20",x"91",x"E3",x"A0",x"01",x"91",x"02",x"29"
		,x"1F",x"C9",x"05",x"F0",x"06",x"A2",x"00",x"8A"
		,x"4C",x"82",x"E8",x"A2",x"00",x"A9",x"01",x"4C"
		,x"82",x"E8",x"20",x"C6",x"E7",x"20",x"A2",x"E3"
		,x"C9",x"FF",x"F0",x"07",x"A2",x"00",x"A9",x"FF"
		,x"4C",x"8C",x"E8",x"A0",x"06",x"B1",x"02",x"8D"
		,x"00",x"B5",x"AD",x"01",x"B5",x"29",x"01",x"D0"
		,x"F9",x"A0",x"05",x"20",x"49",x"E9",x"20",x"28"
		,x"EA",x"A2",x"00",x"86",x"04",x"86",x"05",x"A9"
		,x"18",x"20",x"17",x"EB",x"8D",x"00",x"B5",x"AD"
		,x"01",x"B5",x"29",x"01",x"D0",x"F9",x"A0",x"05"
		,x"20",x"49",x"E9",x"A5",x"04",x"8D",x"00",x"B5"
		,x"AD",x"01",x"B5",x"29",x"01",x"D0",x"F9",x"A0"
		,x"05",x"20",x"49",x"E9",x"8A",x"8D",x"00",x"B5"
		,x"AD",x"01",x"B5",x"29",x"01",x"D0",x"F9",x"A0"
		,x"02",x"B1",x"02",x"8D",x"00",x"B5",x"AD",x"01"
		,x"B5",x"29",x"01",x"D0",x"F9",x"A9",x"95",x"8D"
		,x"00",x"B5",x"AD",x"01",x"B5",x"29",x"01",x"D0"
		,x"F9",x"A0",x"06",x"B1",x"02",x"C9",x"4C",x"D0"
		,x"03",x"20",x"91",x"E3",x"A9",x"0A",x"A0",x"01"
		,x"91",x"02",x"20",x"91",x"E3",x"A0",x"00",x"91"
		,x"02",x"29",x"80",x"F0",x"0B",x"C8",x"38",x"B1"
		,x"02",x"E9",x"01",x"91",x"02",x"AA",x"D0",x"EA"
		,x"A8",x"AA",x"B1",x"02",x"4C",x"8C",x"E8",x"85"
		,x"12",x"A0",x"00",x"B1",x"02",x"85",x"0C",x"85"
		,x"0E",x"C8",x"B1",x"02",x"85",x"0D",x"85",x"0F"
		,x"C8",x"B1",x"02",x"85",x"04",x"C8",x"B1",x"02"
		,x"85",x"05",x"4C",x"36",x"E7",x"20",x"AF",x"E5"
		,x"A4",x"12",x"C0",x"0A",x"D0",x"3C",x"C9",x"00"
		,x"D0",x"11",x"E0",x"80",x"D0",x"0D",x"A0",x"06"
		,x"B9",x"C2",x"F3",x"91",x"0C",x"88",x"10",x"F8"
		,x"4C",x"3E",x"E6",x"A5",x"05",x"10",x"23",x"A9"
		,x"2D",x"A0",x"00",x"91",x"0C",x"E6",x"0C",x"D0"
		,x"02",x"E6",x"0D",x"A5",x"04",x"49",x"FF",x"18"
		,x"69",x"01",x"85",x"04",x"A5",x"05",x"49",x"FF"
		,x"69",x"00",x"85",x"05",x"4C",x"12",x"E6",x"20"
		,x"AF",x"E5",x"A9",x"00",x"48",x"A0",x"10",x"A9"
		,x"00",x"06",x"04",x"26",x"05",x"2A",x"C5",x"12"
		,x"90",x"04",x"E5",x"12",x"E6",x"04",x"88",x"D0"
		,x"F0",x"A8",x"B9",x"B2",x"F3",x"48",x"A5",x"04"
		,x"05",x"05",x"D0",x"E1",x"A0",x"00",x"68",x"91"
		,x"0C",x"F0",x"03",x"C8",x"D0",x"F8",x"A5",x"0E"
		,x"A6",x"0F",x"60",x"49",x"FF",x"85",x"0E",x"8A"
		,x"49",x"FF",x"85",x"0F",x"20",x"62",x"E8",x"85"
		,x"0C",x"86",x"0D",x"20",x"62",x"E8",x"85",x"0A"
		,x"86",x"0B",x"A6",x"0E",x"A0",x"00",x"E8",x"F0"
		,x"0F",x"B1",x"0A",x"D1",x"0C",x"D0",x"10",x"C8"
		,x"D0",x"F4",x"E6",x"0B",x"E6",x"0D",x"D0",x"EE"
		,x"E6",x"0F",x"D0",x"ED",x"4C",x"03",x"ED",x"B0"
		,x"03",x"A2",x"FF",x"60",x"A2",x"01",x"60",x"20"
		,x"9F",x"E6",x"A0",x"00",x"A6",x"0E",x"E8",x"F0"
		,x"0D",x"B1",x"0A",x"91",x"0C",x"C8",x"D0",x"F6"
		,x"E6",x"0B",x"E6",x"0D",x"D0",x"F0",x"E6",x"0F"
		,x"D0",x"EF",x"A5",x"0C",x"A6",x"12",x"60",x"49"
		,x"FF",x"85",x"0E",x"8A",x"49",x"FF",x"85",x"0F"
		,x"20",x"62",x"E8",x"85",x"0A",x"86",x"0B",x"20"
		,x"62",x"E8",x"85",x"0C",x"86",x"0D",x"86",x"12"
		,x"60",x"85",x"0E",x"86",x"0F",x"A9",x"00",x"F0"
		,x"07",x"85",x"0E",x"86",x"0F",x"20",x"62",x"E8"
		,x"85",x"12",x"A0",x"01",x"B1",x"02",x"AA",x"88"
		,x"B1",x"02",x"85",x"0A",x"86",x"0B",x"A5",x"12"
		,x"A0",x"00",x"A6",x"0F",x"F0",x"0D",x"91",x"0A"
		,x"C8",x"91",x"0A",x"C8",x"D0",x"F8",x"E6",x"0B"
		,x"CA",x"D0",x"F3",x"A6",x"0E",x"F0",x"06",x"91"
		,x"0A",x"C8",x"CA",x"D0",x"FA",x"4C",x"62",x"E8"
		,x"A9",x"08",x"85",x"0A",x"A9",x"A0",x"85",x"0B"
		,x"A9",x"00",x"A8",x"A2",x"04",x"F0",x"0A",x"91"
		,x"0A",x"C8",x"D0",x"FB",x"E6",x"0B",x"CA",x"D0"
		,x"F6",x"C0",x"3D",x"F0",x"05",x"91",x"0A",x"C8"
		,x"D0",x"F7",x"60",x"60",x"A2",x"00",x"18",x"A0"
		,x"00",x"71",x"02",x"C8",x"48",x"8A",x"71",x"02"
		,x"AA",x"18",x"A5",x"02",x"69",x"02",x"85",x"02"
		,x"90",x"02",x"E6",x"03",x"68",x"60",x"C8",x"48"
		,x"18",x"98",x"65",x"02",x"85",x"02",x"90",x"02"
		,x"E6",x"03",x"68",x"60",x"A2",x"00",x"A0",x"00"
		,x"31",x"02",x"C8",x"48",x"8A",x"31",x"02",x"AA"
		,x"68",x"4C",x"36",x"E7",x"86",x"12",x"0A",x"26"
		,x"12",x"A6",x"12",x"60",x"86",x"12",x"0A",x"26"
		,x"12",x"0A",x"26",x"12",x"A6",x"12",x"60",x"86"
		,x"12",x"0A",x"26",x"12",x"0A",x"26",x"12",x"0A"
		,x"26",x"12",x"A6",x"12",x"60",x"85",x"0A",x"86"
		,x"0B",x"6C",x"0A",x"00",x"49",x"FF",x"48",x"8A"
		,x"49",x"FF",x"AA",x"68",x"60",x"A9",x"C9",x"A2"
		,x"F3",x"A0",x"00",x"D0",x"0A",x"60",x"A9",x"C9"
		,x"A2",x"F3",x"A0",x"00",x"D0",x"01",x"60",x"8D"
		,x"02",x"A0",x"8E",x"03",x"A0",x"8C",x"44",x"A4"
		,x"AC",x"44",x"A4",x"F0",x"17",x"88",x"20",x"01"
		,x"A0",x"8D",x"07",x"A0",x"88",x"20",x"01",x"A0"
		,x"8D",x"06",x"A0",x"8C",x"44",x"A4",x"20",x"05"
		,x"A0",x"4C",x"A0",x"E7",x"60",x"A4",x"02",x"D0"
		,x"02",x"C6",x"03",x"C6",x"02",x"60",x"A5",x"02"
		,x"38",x"E9",x"02",x"85",x"02",x"90",x"01",x"60"
		,x"C6",x"03",x"60",x"A5",x"02",x"38",x"E9",x"03"
		,x"85",x"02",x"90",x"01",x"60",x"C6",x"03",x"60"
		,x"A5",x"02",x"38",x"E9",x"04",x"85",x"02",x"90"
		,x"01",x"60",x"C6",x"03",x"60",x"A5",x"02",x"38"
		,x"E9",x"05",x"85",x"02",x"90",x"01",x"60",x"C6"
		,x"03",x"60",x"A5",x"02",x"38",x"E9",x"06",x"85"
		,x"02",x"90",x"01",x"60",x"C6",x"03",x"60",x"A5"
		,x"02",x"38",x"E9",x"07",x"85",x"02",x"90",x"01"
		,x"60",x"C6",x"03",x"60",x"A5",x"02",x"38",x"E9"
		,x"08",x"85",x"02",x"90",x"01",x"60",x"C6",x"03"
		,x"60",x"98",x"A4",x"02",x"D0",x"02",x"C6",x"03"
		,x"C6",x"02",x"A0",x"00",x"91",x"02",x"60",x"85"
		,x"04",x"86",x"05",x"A0",x"00",x"B1",x"02",x"AA"
		,x"E6",x"02",x"D0",x"02",x"E6",x"03",x"B1",x"02"
		,x"E6",x"02",x"D0",x"02",x"E6",x"03",x"38",x"E5"
		,x"05",x"D0",x"09",x"E4",x"04",x"F0",x"04",x"69"
		,x"FF",x"09",x"01",x"60",x"50",x"FD",x"49",x"FF"
		,x"09",x"01",x"60",x"E6",x"02",x"D0",x"02",x"E6"
		,x"03",x"60",x"A0",x"01",x"B1",x"02",x"AA",x"88"
		,x"B1",x"02",x"E6",x"02",x"F0",x"05",x"E6",x"02"
		,x"F0",x"03",x"60",x"E6",x"02",x"E6",x"03",x"60"
		,x"A0",x"03",x"4C",x"37",x"E7",x"A0",x"04",x"4C"
		,x"37",x"E7",x"A0",x"05",x"4C",x"37",x"E7",x"A0"
		,x"06",x"4C",x"37",x"E7",x"A0",x"07",x"4C",x"37"
		,x"E7",x"A0",x"00",x"18",x"71",x"02",x"85",x"12"
		,x"C8",x"8A",x"71",x"02",x"AA",x"C8",x"A5",x"04"
		,x"71",x"02",x"85",x"04",x"C8",x"A5",x"05",x"71"
		,x"02",x"85",x"05",x"A5",x"12",x"4C",x"36",x"E7"
		,x"A0",x"00",x"31",x"02",x"85",x"12",x"C8",x"8A"
		,x"31",x"02",x"AA",x"C8",x"A5",x"04",x"31",x"02"
		,x"85",x"04",x"C8",x"A5",x"05",x"31",x"02",x"85"
		,x"05",x"A5",x"12",x"4C",x"36",x"E7",x"86",x"12"
		,x"A2",x"00",x"05",x"12",x"05",x"04",x"05",x"05"
		,x"D0",x"03",x"A9",x"01",x"60",x"8A",x"60",x"85"
		,x"0A",x"86",x"0B",x"A0",x"03",x"B1",x"02",x"38"
		,x"E5",x"05",x"D0",x"22",x"88",x"B1",x"02",x"C5"
		,x"04",x"D0",x"0C",x"88",x"B1",x"02",x"C5",x"0B"
		,x"D0",x"05",x"88",x"B1",x"02",x"C5",x"0A",x"08"
		,x"20",x"7D",x"E8",x"28",x"F0",x"04",x"B0",x"03"
		,x"A9",x"FF",x"60",x"A9",x"01",x"60",x"50",x"04"
		,x"49",x"FF",x"09",x"01",x"08",x"20",x"7D",x"E8"
		,x"28",x"60",x"A0",x"01",x"85",x"0A",x"86",x"0B"
		,x"B1",x"0A",x"AA",x"88",x"B1",x"0A",x"60",x"A0"
		,x"01",x"B1",x"02",x"AA",x"88",x"B1",x"02",x"60"
		,x"A0",x"03",x"85",x"0A",x"86",x"0B",x"B1",x"0A"
		,x"88",x"85",x"05",x"B1",x"0A",x"88",x"85",x"04"
		,x"B1",x"0A",x"88",x"AA",x"B1",x"0A",x"60",x"A0"
		,x"03",x"B1",x"02",x"85",x"05",x"88",x"B1",x"02"
		,x"85",x"04",x"88",x"B1",x"02",x"AA",x"88",x"B1"
		,x"02",x"60",x"84",x"12",x"38",x"E5",x"12",x"85"
		,x"12",x"8A",x"E9",x"00",x"AA",x"A5",x"04",x"E9"
		,x"00",x"85",x"04",x"A5",x"05",x"E9",x"00",x"85"
		,x"05",x"A5",x"12",x"60",x"A9",x"00",x"A2",x"00"
		,x"F0",x"07",x"A9",x"00",x"A2",x"00",x"20",x"37"
		,x"E7",x"48",x"A0",x"00",x"B1",x"02",x"38",x"65"
		,x"02",x"85",x"02",x"90",x"02",x"E6",x"03",x"68"
		,x"60",x"20",x"DF",x"E8",x"4C",x"6B",x"EC",x"84"
		,x"10",x"18",x"65",x"10",x"90",x"09",x"E8",x"D0"
		,x"06",x"E6",x"04",x"D0",x"02",x"E6",x"05",x"60"
		,x"85",x"0A",x"86",x"0B",x"A0",x"00",x"B1",x"02"
		,x"85",x"0E",x"C8",x"B1",x"02",x"85",x"0F",x"C8"
		,x"B1",x"02",x"85",x"10",x"C8",x"B1",x"02",x"85"
		,x"11",x"20",x"36",x"E7",x"A9",x"00",x"85",x"15"
		,x"85",x"14",x"85",x"13",x"A0",x"20",x"46",x"15"
		,x"66",x"14",x"66",x"13",x"6A",x"66",x"05",x"66"
		,x"04",x"66",x"0B",x"66",x"0A",x"90",x"17",x"18"
		,x"65",x"0E",x"48",x"A5",x"0F",x"65",x"13",x"85"
		,x"13",x"A5",x"10",x"65",x"14",x"85",x"14",x"A5"
		,x"11",x"65",x"15",x"85",x"15",x"68",x"88",x"10"
		,x"D5",x"A5",x"0A",x"A6",x"0B",x"60",x"20",x"DF"
		,x"E8",x"4C",x"65",x"EC",x"A0",x"00",x"11",x"02"
		,x"85",x"12",x"C8",x"8A",x"11",x"02",x"AA",x"C8"
		,x"A5",x"04",x"11",x"02",x"85",x"04",x"C8",x"A5"
		,x"05",x"11",x"02",x"85",x"05",x"A5",x"12",x"4C"
		,x"36",x"E7",x"A0",x"00",x"84",x"04",x"84",x"05"
		,x"48",x"20",x"E0",x"E7",x"A0",x"03",x"A5",x"05"
		,x"91",x"02",x"88",x"A5",x"04",x"91",x"02",x"88"
		,x"8A",x"91",x"02",x"88",x"68",x"91",x"02",x"60"
		,x"85",x"06",x"86",x"07",x"A5",x"04",x"85",x"08"
		,x"A5",x"05",x"85",x"09",x"A5",x"06",x"60",x"A5"
		,x"09",x"85",x"05",x"A5",x"08",x"85",x"04",x"A6"
		,x"07",x"A5",x"06",x"60",x"48",x"A0",x"00",x"B1"
		,x"02",x"85",x"0A",x"C8",x"B1",x"02",x"85",x"0B"
		,x"C8",x"B1",x"02",x"85",x"0C",x"C8",x"B1",x"02"
		,x"85",x"0D",x"68",x"20",x"36",x"E7",x"A8",x"8A"
		,x"05",x"04",x"05",x"05",x"D0",x"3D",x"C0",x"20"
		,x"B0",x"39",x"C0",x"00",x"F0",x"34",x"98",x"C9"
		,x"08",x"90",x"14",x"E9",x"08",x"A6",x"0C",x"86"
		,x"0D",x"A6",x"0B",x"86",x"0C",x"A6",x"0A",x"86"
		,x"0B",x"A2",x"00",x"86",x"0A",x"F0",x"E8",x"A8"
		,x"A5",x"0A",x"C0",x"00",x"F0",x"0A",x"0A",x"26"
		,x"0B",x"26",x"0C",x"26",x"0D",x"88",x"D0",x"F6"
		,x"A6",x"0C",x"86",x"04",x"A6",x"0D",x"86",x"05"
		,x"A6",x"0B",x"60",x"A9",x"00",x"85",x"05",x"85"
		,x"04",x"AA",x"60",x"20",x"60",x"EB",x"20",x"7A"
		,x"EB",x"B0",x"3F",x"C0",x"00",x"F0",x"3A",x"98"
		,x"C9",x"08",x"90",x"18",x"E9",x"08",x"A6",x"0B"
		,x"86",x"0A",x"A6",x"0C",x"86",x"0B",x"A0",x"00"
		,x"A6",x"0D",x"86",x"0C",x"10",x"01",x"88",x"84"
		,x"0D",x"4C",x"D0",x"EA",x"A8",x"A5",x"0D",x"C0"
		,x"00",x"F0",x"0C",x"C9",x"80",x"6A",x"66",x"0C"
		,x"66",x"0B",x"66",x"0A",x"88",x"D0",x"F4",x"85"
		,x"05",x"A5",x"0C",x"85",x"04",x"A6",x"0B",x"A5"
		,x"0A",x"60",x"A2",x"00",x"A5",x"0D",x"10",x"01"
		,x"CA",x"86",x"05",x"86",x"04",x"8A",x"60",x"20"
		,x"60",x"EB",x"20",x"7A",x"EB",x"B0",x"39",x"C0"
		,x"00",x"F0",x"34",x"98",x"C9",x"08",x"90",x"14"
		,x"E9",x"08",x"A6",x"0B",x"86",x"0A",x"A6",x"0C"
		,x"86",x"0B",x"A6",x"0D",x"86",x"0C",x"A2",x"00"
		,x"86",x"0D",x"F0",x"E8",x"A8",x"A5",x"0D",x"C0"
		,x"00",x"F0",x"0A",x"4A",x"66",x"0C",x"66",x"0B"
		,x"66",x"0A",x"88",x"D0",x"F6",x"85",x"05",x"A5"
		,x"0C",x"85",x"04",x"A6",x"0B",x"A5",x"0A",x"60"
		,x"A9",x"00",x"85",x"05",x"85",x"04",x"AA",x"60"
		,x"48",x"A0",x"00",x"B1",x"02",x"85",x"0A",x"C8"
		,x"B1",x"02",x"85",x"0B",x"C8",x"B1",x"02",x"85"
		,x"0C",x"C8",x"B1",x"02",x"85",x"0D",x"68",x"4C"
		,x"36",x"E7",x"A8",x"8A",x"05",x"04",x"05",x"05"
		,x"D0",x"04",x"C0",x"20",x"90",x"01",x"38",x"60"
		,x"A0",x"00",x"38",x"49",x"FF",x"71",x"02",x"91"
		,x"02",x"48",x"C8",x"8A",x"49",x"FF",x"71",x"02"
		,x"91",x"02",x"AA",x"C8",x"B1",x"02",x"E5",x"04"
		,x"91",x"02",x"85",x"04",x"C8",x"B1",x"02",x"E5"
		,x"05",x"91",x"02",x"85",x"05",x"68",x"60",x"A0"
		,x"00",x"38",x"49",x"FF",x"71",x"02",x"48",x"C8"
		,x"8A",x"49",x"FF",x"71",x"02",x"AA",x"C8",x"B1"
		,x"02",x"E5",x"04",x"85",x"04",x"C8",x"B1",x"02"
		,x"E5",x"05",x"85",x"05",x"68",x"4C",x"36",x"E7"
		,x"A8",x"86",x"12",x"05",x"12",x"05",x"04",x"05"
		,x"05",x"F0",x"03",x"98",x"A0",x"01",x"60",x"20"
		,x"EA",x"EB",x"20",x"0E",x"EC",x"A5",x"0A",x"A6"
		,x"0B",x"60",x"85",x"0E",x"86",x"0F",x"A5",x"04"
		,x"85",x"10",x"A5",x"05",x"85",x"11",x"A0",x"00"
		,x"B1",x"02",x"85",x"0A",x"C8",x"B1",x"02",x"85"
		,x"0B",x"C8",x"B1",x"02",x"85",x"04",x"C8",x"B1"
		,x"02",x"85",x"05",x"4C",x"36",x"E7",x"A9",x"00"
		,x"85",x"0D",x"85",x"14",x"85",x"15",x"A0",x"20"
		,x"06",x"0A",x"26",x"0B",x"26",x"04",x"26",x"05"
		,x"2A",x"26",x"0D",x"26",x"14",x"26",x"15",x"48"
		,x"C5",x"0E",x"A5",x"0D",x"E5",x"0F",x"A5",x"14"
		,x"E5",x"10",x"A5",x"15",x"E5",x"11",x"90",x"14"
		,x"85",x"11",x"68",x"E5",x"0E",x"48",x"A5",x"0D"
		,x"E5",x"0F",x"85",x"0D",x"A5",x"14",x"E5",x"10"
		,x"85",x"14",x"E6",x"0A",x"68",x"88",x"D0",x"C8"
		,x"85",x"0C",x"60",x"20",x"DF",x"E8",x"4C",x"8B"
		,x"EC",x"20",x"DF",x"E8",x"4C",x"89",x"EC",x"20"
		,x"DF",x"E8",x"4C",x"83",x"EC",x"D0",x"2A",x"A2"
		,x"00",x"8A",x"60",x"F0",x"24",x"A2",x"00",x"8A"
		,x"60",x"F0",x"1E",x"30",x"1C",x"A2",x"00",x"8A"
		,x"60",x"F0",x"02",x"10",x"14",x"A2",x"00",x"8A"
		,x"60",x"F0",x"0E",x"90",x"0C",x"A2",x"00",x"8A"
		,x"60",x"F0",x"02",x"B0",x"04",x"A2",x"00",x"8A"
		,x"60",x"A2",x"00",x"A9",x"01",x"60",x"85",x"0A"
		,x"86",x"0B",x"0A",x"26",x"0B",x"18",x"65",x"0A"
		,x"48",x"8A",x"65",x"0B",x"AA",x"68",x"60",x"48"
		,x"A0",x"00",x"B1",x"02",x"85",x"04",x"C8",x"B1"
		,x"02",x"85",x"05",x"68",x"4C",x"6A",x"E8",x"A0"
		,x"00",x"B1",x"02",x"A4",x"02",x"F0",x"07",x"C6"
		,x"02",x"A0",x"00",x"91",x"02",x"60",x"C6",x"03"
		,x"C6",x"02",x"91",x"02",x"60",x"A9",x"00",x"A2"
		,x"00",x"48",x"A5",x"02",x"38",x"E9",x"02",x"85"
		,x"02",x"B0",x"02",x"C6",x"03",x"A0",x"01",x"8A"
		,x"91",x"02",x"68",x"88",x"91",x"02",x"60",x"A0"
		,x"03",x"A5",x"02",x"38",x"E9",x"02",x"85",x"02"
		,x"B0",x"02",x"C6",x"03",x"B1",x"02",x"AA",x"88"
		,x"B1",x"02",x"A0",x"00",x"91",x"02",x"C8",x"8A"
		,x"91",x"02",x"60",x"A9",x"00",x"AA",x"60",x"A2"
		,x"00",x"20",x"A7",x"EC",x"E0",x"00",x"D0",x"2A"
		,x"C9",x"10",x"B0",x"26",x"C9",x"08",x"F0",x"19"
		,x"90",x"09",x"A4",x"04",x"84",x"05",x"86",x"04"
		,x"38",x"E9",x"08",x"A8",x"F0",x"0F",x"A5",x"04"
		,x"0A",x"26",x"05",x"88",x"D0",x"FA",x"A6",x"05"
		,x"60",x"8A",x"A6",x"04",x"60",x"A5",x"04",x"A6"
		,x"05",x"60",x"4C",x"03",x"ED",x"86",x"12",x"46"
		,x"12",x"6A",x"A6",x"12",x"60",x"86",x"12",x"46"
		,x"12",x"6A",x"46",x"12",x"6A",x"46",x"12",x"6A"
		,x"46",x"12",x"6A",x"A6",x"12",x"60",x"A2",x"00"
		,x"20",x"A7",x"EC",x"E0",x"00",x"D0",x"35",x"C9"
		,x"10",x"B0",x"31",x"C9",x"08",x"F0",x"22",x"90"
		,x"0E",x"A0",x"00",x"A6",x"05",x"86",x"04",x"10"
		,x"01",x"88",x"84",x"05",x"38",x"E9",x"08",x"A8"
		,x"F0",x"15",x"A5",x"04",x"A6",x"05",x"E0",x"80"
		,x"66",x"05",x"6A",x"88",x"D0",x"F8",x"A6",x"05"
		,x"60",x"A5",x"05",x"10",x"01",x"CA",x"60",x"A5"
		,x"04",x"A6",x"05",x"60",x"4C",x"03",x"ED",x"A2"
		,x"00",x"20",x"A7",x"EC",x"E0",x"00",x"D0",x"F4"
		,x"C9",x"10",x"B0",x"F0",x"C9",x"08",x"F0",x"18"
		,x"90",x"08",x"E9",x"08",x"A4",x"05",x"84",x"04"
		,x"86",x"05",x"A8",x"F0",x"DA",x"A5",x"04",x"46"
		,x"05",x"6A",x"88",x"D0",x"FA",x"A6",x"05",x"60"
		,x"A5",x"05",x"60",x"48",x"84",x"12",x"A0",x"01"
		,x"B1",x"02",x"85",x"0B",x"88",x"B1",x"02",x"85"
		,x"0A",x"A4",x"12",x"68",x"91",x"0A",x"4C",x"6A"
		,x"E8",x"A0",x"00",x"91",x"02",x"C8",x"48",x"8A"
		,x"91",x"02",x"68",x"60",x"85",x"12",x"86",x"13"
		,x"84",x"14",x"20",x"62",x"E8",x"85",x"0A",x"86"
		,x"0B",x"A4",x"14",x"A5",x"12",x"91",x"0A",x"C8"
		,x"A5",x"13",x"91",x"0A",x"C8",x"AA",x"A5",x"04"
		,x"91",x"0A",x"C8",x"A5",x"05",x"91",x"0A",x"A5"
		,x"12",x"60",x"A0",x"00",x"91",x"02",x"C8",x"48"
		,x"8A",x"91",x"02",x"C8",x"A5",x"04",x"91",x"02"
		,x"C8",x"A5",x"05",x"91",x"02",x"68",x"60",x"A0"
		,x"00",x"38",x"49",x"FF",x"71",x"02",x"91",x"02"
		,x"48",x"C8",x"8A",x"49",x"FF",x"71",x"02",x"91"
		,x"02",x"AA",x"68",x"60",x"A2",x"00",x"38",x"49"
		,x"FF",x"A0",x"00",x"71",x"02",x"C8",x"48",x"8A"
		,x"49",x"FF",x"71",x"02",x"AA",x"68",x"4C",x"36"
		,x"E7",x"98",x"49",x"FF",x"38",x"65",x"02",x"85"
		,x"02",x"B0",x"02",x"C6",x"03",x"60",x"48",x"20"
		,x"C6",x"E7",x"A0",x"02",x"B1",x"02",x"A0",x"00"
		,x"91",x"02",x"A0",x"03",x"B1",x"02",x"A0",x"01"
		,x"91",x"02",x"A9",x"00",x"C8",x"91",x"02",x"C8"
		,x"91",x"02",x"68",x"60",x"48",x"20",x"C6",x"E7"
		,x"A0",x"02",x"B1",x"02",x"A0",x"00",x"91",x"02"
		,x"A0",x"03",x"B1",x"02",x"10",x"E0",x"A0",x"01"
		,x"91",x"02",x"A9",x"FF",x"D0",x"DE",x"A2",x"00"
		,x"85",x"10",x"86",x"11",x"20",x"A7",x"EC",x"20"
		,x"9F",x"EE",x"A5",x"04",x"A6",x"05",x"60",x"A9"
		,x"00",x"85",x"0B",x"A0",x"10",x"06",x"04",x"26"
		,x"05",x"2A",x"26",x"0B",x"48",x"C5",x"10",x"A5"
		,x"0B",x"E5",x"11",x"90",x"08",x"85",x"0B",x"68"
		,x"E5",x"10",x"48",x"E6",x"04",x"68",x"88",x"D0"
		,x"E4",x"85",x"0A",x"60",x"A2",x"00",x"85",x"10"
		,x"86",x"11",x"20",x"A7",x"EC",x"20",x"9F",x"EE"
		,x"A5",x"0A",x"A6",x"0B",x"60",x"42",x"6F",x"6F"
		,x"74",x"6C",x"6F",x"61",x"64",x"65",x"72",x"3E"
		,x"0A",x"0D",x"00",x"2A",x"20",x"46",x"50",x"47"
		,x"41",x"20",x"46",x"6C",x"6F",x"70",x"70",x"79"
		,x"20",x"20",x"2A",x"0A",x"62",x"6F",x"6F",x"74"
		,x"69",x"6E",x"67",x"2E",x"2E",x"2E",x"0A",x"00"
		,x"73",x"77",x"69",x"74",x"63",x"68",x"20",x"36"
		,x"20",x"6F",x"6E",x"20",x"2D",x"0A",x"00",x"49"
		,x"6E",x"69",x"74",x"69",x"6E",x"67",x"20",x"4D"
		,x"4D",x"43",x"2E",x"2E",x"2E",x"0A",x"00",x"73"
		,x"79",x"73",x"2F",x"66",x"69",x"72",x"6D",x"77"
		,x"61",x"72",x"65",x"2E",x"62",x"69",x"6E",x"00"
		,x"73",x"79",x"73",x"2F",x"66",x"69",x"72",x"6D"
		,x"77",x"61",x"72",x"65",x"2E",x"62",x"69",x"6E"
		,x"0A",x"6E",x"6F",x"74",x"20",x"66",x"6F",x"75"
		,x"6E",x"64",x"2E",x"0A",x"00",x"6E",x"6F",x"20"
		,x"4D",x"4D",x"43",x"2F",x"53",x"44",x"20",x"63"
		,x"61",x"72",x"64",x"2E",x"0A",x"00",x"6E",x"6F"
		,x"20",x"46",x"41",x"54",x"0A",x"66",x"69",x"6C"
		,x"65",x"73",x"79",x"73",x"74",x"65",x"6D",x"2E"
		,x"0A",x"00",x"4C",x"6F",x"61",x"64",x"69",x"6E"
		,x"67",x"0A",x"66",x"69",x"72",x"6D",x"77",x"61"
		,x"72",x"65",x"2E",x"2E",x"2E",x"0A",x"00",x"55"
		,x"61",x"72",x"74",x"20",x"6D",x"6F",x"64",x"65"
		,x"2E",x"00",x"52",x"45",x"41",x"44",x"59",x"2E"
		,x"0D",x"0A",x"00",x"30",x"00",x"20",x"00",x"0D"
		,x"0A",x"00",x"46",x"41",x"54",x"31",x"32",x"46"
		,x"41",x"54",x"31",x"36",x"46",x"41",x"54",x"33"
		,x"32",x"00",x"00",x"3E",x"7F",x"41",x"4D",x"4F"
		,x"2E",x"00",x"00",x"20",x"74",x"54",x"54",x"7C"
		,x"78",x"00",x"00",x"7E",x"7E",x"48",x"48",x"78"
		,x"30",x"00",x"00",x"38",x"7C",x"44",x"44",x"44"
		,x"00",x"00",x"00",x"30",x"78",x"48",x"48",x"7E"
		,x"7E",x"00",x"00",x"38",x"7C",x"54",x"54",x"5C"
		,x"18",x"00",x"00",x"00",x"08",x"7C",x"7E",x"0A"
		,x"0A",x"00",x"00",x"98",x"BC",x"A4",x"A4",x"FC"
		,x"7C",x"00",x"00",x"7E",x"7E",x"08",x"08",x"78"
		,x"70",x"00",x"00",x"00",x"48",x"7A",x"7A",x"40"
		,x"00",x"00",x"00",x"00",x"80",x"80",x"80",x"FA"
		,x"7A",x"00",x"00",x"7E",x"7E",x"10",x"38",x"68"
		,x"40",x"00",x"00",x"00",x"42",x"7E",x"7E",x"40"
		,x"00",x"00",x"00",x"7C",x"7C",x"18",x"38",x"1C"
		,x"7C",x"78",x"00",x"7C",x"7C",x"04",x"04",x"7C"
		,x"78",x"00",x"00",x"38",x"7C",x"44",x"44",x"7C"
		,x"38",x"00",x"00",x"FC",x"FC",x"24",x"24",x"3C"
		,x"18",x"00",x"00",x"18",x"3C",x"24",x"24",x"FC"
		,x"FC",x"00",x"00",x"7C",x"7C",x"04",x"04",x"0C"
		,x"08",x"00",x"00",x"48",x"5C",x"54",x"54",x"74"
		,x"24",x"00",x"00",x"04",x"04",x"3E",x"7E",x"44"
		,x"44",x"00",x"00",x"3C",x"7C",x"40",x"40",x"7C"
		,x"7C",x"00",x"00",x"1C",x"3C",x"60",x"60",x"3C"
		,x"1C",x"00",x"00",x"1C",x"7C",x"70",x"38",x"70"
		,x"7C",x"1C",x"00",x"44",x"6C",x"38",x"38",x"6C"
		,x"44",x"00",x"00",x"9C",x"BC",x"A0",x"E0",x"7C"
		,x"3C",x"00",x"00",x"44",x"64",x"74",x"5C",x"4C"
		,x"44",x"00",x"00",x"00",x"7F",x"7F",x"41",x"41"
		,x"00",x"00",x"40",x"68",x"7C",x"5E",x"49",x"49"
		,x"22",x"00",x"00",x"00",x"41",x"41",x"7F",x"7F"
		,x"00",x"00",x"00",x"08",x"0C",x"FE",x"FE",x"0C"
		,x"08",x"00",x"00",x"18",x"3C",x"7E",x"18",x"18"
		,x"18",x"18",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"4F",x"4F",x"00"
		,x"00",x"00",x"00",x"07",x"07",x"00",x"00",x"07"
		,x"07",x"00",x"14",x"7F",x"7F",x"14",x"14",x"7F"
		,x"7F",x"14",x"00",x"24",x"2E",x"6B",x"6B",x"3A"
		,x"12",x"00",x"00",x"63",x"33",x"18",x"0C",x"66"
		,x"63",x"00",x"00",x"32",x"7F",x"4D",x"4D",x"77"
		,x"72",x"50",x"00",x"00",x"00",x"04",x"06",x"03"
		,x"01",x"00",x"00",x"00",x"1C",x"3E",x"63",x"41"
		,x"00",x"00",x"00",x"00",x"41",x"63",x"3E",x"1C"
		,x"00",x"00",x"08",x"2A",x"3E",x"1C",x"1C",x"3E"
		,x"2A",x"08",x"00",x"08",x"08",x"3E",x"3E",x"08"
		,x"08",x"00",x"00",x"00",x"80",x"E0",x"60",x"00"
		,x"00",x"00",x"00",x"08",x"08",x"08",x"08",x"08"
		,x"08",x"00",x"00",x"00",x"00",x"60",x"60",x"00"
		,x"00",x"00",x"00",x"40",x"60",x"30",x"18",x"0C"
		,x"06",x"02",x"00",x"3E",x"7F",x"49",x"45",x"7F"
		,x"3E",x"00",x"00",x"40",x"44",x"7F",x"7F",x"40"
		,x"40",x"00",x"00",x"62",x"73",x"51",x"49",x"4F"
		,x"46",x"00",x"00",x"22",x"63",x"49",x"49",x"7F"
		,x"36",x"00",x"00",x"18",x"18",x"14",x"16",x"7F"
		,x"7F",x"10",x"00",x"27",x"67",x"45",x"45",x"7D"
		,x"39",x"00",x"00",x"3E",x"7F",x"49",x"49",x"7B"
		,x"32",x"00",x"00",x"03",x"03",x"79",x"7D",x"07"
		,x"03",x"00",x"00",x"36",x"7F",x"49",x"49",x"7F"
		,x"36",x"00",x"00",x"26",x"6F",x"49",x"49",x"7F"
		,x"3E",x"00",x"00",x"00",x"00",x"24",x"24",x"00"
		,x"00",x"00",x"00",x"00",x"80",x"E4",x"64",x"00"
		,x"00",x"00",x"00",x"08",x"1C",x"36",x"63",x"41"
		,x"41",x"00",x"00",x"14",x"14",x"14",x"14",x"14"
		,x"14",x"00",x"00",x"41",x"41",x"63",x"36",x"1C"
		,x"08",x"00",x"00",x"02",x"03",x"51",x"59",x"0F"
		,x"06",x"00",x"18",x"18",x"18",x"18",x"18",x"18"
		,x"18",x"18",x"00",x"7C",x"7E",x"0B",x"0B",x"7E"
		,x"7C",x"00",x"00",x"7F",x"7F",x"49",x"49",x"7F"
		,x"36",x"00",x"00",x"3E",x"7F",x"41",x"41",x"63"
		,x"22",x"00",x"00",x"7F",x"7F",x"41",x"63",x"3E"
		,x"1C",x"00",x"00",x"7F",x"7F",x"49",x"49",x"41"
		,x"41",x"00",x"00",x"7F",x"7F",x"09",x"09",x"01"
		,x"01",x"00",x"00",x"3E",x"7F",x"41",x"49",x"7B"
		,x"3A",x"00",x"00",x"7F",x"7F",x"08",x"08",x"7F"
		,x"7F",x"00",x"00",x"00",x"41",x"7F",x"7F",x"41"
		,x"00",x"00",x"00",x"20",x"60",x"41",x"7F",x"3F"
		,x"01",x"00",x"00",x"7F",x"7F",x"1C",x"36",x"63"
		,x"41",x"00",x"00",x"7F",x"7F",x"40",x"40",x"40"
		,x"40",x"00",x"00",x"7F",x"7F",x"06",x"0C",x"06"
		,x"7F",x"7F",x"00",x"7F",x"7F",x"0E",x"1C",x"7F"
		,x"7F",x"00",x"00",x"3E",x"7F",x"41",x"41",x"7F"
		,x"3E",x"00",x"00",x"7F",x"7F",x"09",x"09",x"0F"
		,x"06",x"00",x"00",x"1E",x"3F",x"21",x"61",x"7F"
		,x"5E",x"00",x"00",x"7F",x"7F",x"19",x"39",x"6F"
		,x"46",x"00",x"00",x"26",x"6F",x"49",x"49",x"7B"
		,x"32",x"00",x"00",x"01",x"01",x"7F",x"7F",x"01"
		,x"01",x"00",x"00",x"3F",x"7F",x"40",x"40",x"7F"
		,x"3F",x"00",x"00",x"1F",x"3F",x"60",x"60",x"3F"
		,x"1F",x"00",x"00",x"7F",x"7F",x"30",x"18",x"30"
		,x"7F",x"7F",x"00",x"63",x"77",x"1C",x"1C",x"77"
		,x"63",x"00",x"00",x"07",x"0F",x"78",x"78",x"0F"
		,x"07",x"00",x"00",x"61",x"71",x"59",x"4D",x"47"
		,x"43",x"00",x"18",x"18",x"18",x"FF",x"FF",x"18"
		,x"18",x"18",x"33",x"33",x"CC",x"CC",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00"
		,x"00",x"00",x"CC",x"CC",x"33",x"33",x"CC",x"CC"
		,x"33",x"33",x"66",x"CC",x"99",x"33",x"66",x"CC"
		,x"99",x"33",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00"
		,x"00",x"00",x"F0",x"F0",x"F0",x"F0",x"F0",x"F0"
		,x"F0",x"F0",x"01",x"01",x"01",x"01",x"01",x"01"
		,x"01",x"01",x"80",x"80",x"80",x"80",x"80",x"80"
		,x"80",x"80",x"FF",x"FF",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"33",x"33",x"CC",x"CC",x"33",x"33"
		,x"CC",x"CC",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"FF",x"FF",x"30",x"30",x"C0",x"C0",x"30",x"30"
		,x"C0",x"C0",x"33",x"99",x"CC",x"66",x"33",x"99"
		,x"CC",x"66",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"FF",x"FF",x"00",x"00",x"00",x"FF",x"FF",x"18"
		,x"18",x"18",x"00",x"00",x"00",x"00",x"F0",x"F0"
		,x"F0",x"F0",x"00",x"00",x"00",x"1F",x"1F",x"18"
		,x"18",x"18",x"18",x"18",x"18",x"F8",x"F8",x"00"
		,x"00",x"00",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0"
		,x"C0",x"C0",x"00",x"00",x"00",x"F8",x"F8",x"18"
		,x"18",x"18",x"18",x"18",x"18",x"1F",x"1F",x"18"
		,x"18",x"18",x"18",x"18",x"18",x"F8",x"F8",x"18"
		,x"18",x"18",x"18",x"18",x"18",x"FF",x"FF",x"00"
		,x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF"
		,x"FF",x"FF",x"03",x"03",x"03",x"03",x"03",x"03"
		,x"03",x"03",x"07",x"07",x"07",x"07",x"07",x"07"
		,x"07",x"07",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0"
		,x"E0",x"E0",x"00",x"78",x"78",x"30",x"18",x"0C"
		,x"06",x"03",x"F0",x"F0",x"F0",x"F0",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"0F"
		,x"0F",x"0F",x"18",x"18",x"18",x"1F",x"1F",x"00"
		,x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"00",x"00"
		,x"00",x"00",x"0F",x"0F",x"0F",x"0F",x"F0",x"F0"
		,x"F0",x"F0",x"30",x"31",x"32",x"33",x"34",x"35"
		,x"36",x"37",x"38",x"39",x"41",x"42",x"43",x"44"
		,x"45",x"46",x"2D",x"33",x"32",x"37",x"36",x"38"
		,x"00",x"01",x"B9",x"FF",x"FF",x"60",x"4C",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"
		,x"00",x"00",x"00",x"00",x"00",x"C0",x"00",x"C0"
			);
begin
	p_rom : process(clk, addr)
	begin
	if clk'event and clk = '0' then
		data <= ROM(to_integer(unsigned(addr)));
	end if;
	end process;
end rtl;
