
library ieee;
use ieee.std_logic_1164.all;

use ieee.numeric_std.all;

entity rom is
port (addr	:in std_logic_vector (13 downto 0);
        data  :out std_logic_vector (7 downto 0); 
		  clk :in std_logic );
end rom;


architecture rtl of rom is
	type rom_array is array (0 to 16383) of std_logic_vector(7 downto 0);
constant ROM : ROM_ARRAY := (
		x"97",x"E0",x"43",x"4F",x"50",x"59",x"52",x"49"
		,x"47",x"48",x"54",x"20",x"28",x"43",x"29",x"31"
		,x"39",x"38",x"32",x"2C",x"31",x"39",x"38",x"35"
		,x"2C",x"31",x"39",x"38",x"37",x"20",x"43",x"4F"
		,x"4D",x"4D",x"4F",x"44",x"4F",x"52",x"45",x"20"
		,x"45",x"4C",x"45",x"43",x"54",x"52",x"4F",x"4E"
		,x"49",x"43",x"53",x"2C",x"20",x"4C",x"54",x"44"
		,x"2E",x"0D",x"41",x"4C",x"4C",x"20",x"52",x"49"
		,x"47",x"48",x"54",x"53",x"20",x"52",x"45",x"53"
		,x"45",x"52",x"56",x"45",x"44",x"0D",x"AD",x"0C"
		,x"1C",x"29",x"1F",x"09",x"C0",x"8D",x"0C",x"1C"
		,x"A9",x"FF",x"8D",x"03",x"1C",x"A9",x"55",x"8D"
		,x"01",x"1C",x"A2",x"03",x"A0",x"00",x"50",x"FE"
		,x"B8",x"88",x"D0",x"FA",x"CA",x"D0",x"F7",x"60"
		,x"A4",x"82",x"4C",x"EE",x"D3",x"95",x"B5",x"95"
		,x"BB",x"A9",x"00",x"9D",x"44",x"02",x"60",x"08"
		,x"78",x"A9",x"00",x"F8",x"E0",x"00",x"F0",x"07"
		,x"18",x"69",x"01",x"CA",x"4C",x"84",x"C0",x"28"
		,x"4C",x"AA",x"E6",x"C9",x"03",x"B0",x"05",x"A9"
		,x"72",x"20",x"C7",x"E6",x"A9",x"01",x"60",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"78",x"A9",x"F7",x"2D",x"00",x"1C",x"48",x"A5"
		,x"7F",x"F0",x"05",x"68",x"09",x"00",x"D0",x"03"
		,x"68",x"09",x"08",x"8D",x"00",x"1C",x"58",x"60"
		,x"78",x"A9",x"08",x"0D",x"00",x"1C",x"8D",x"00"
		,x"1C",x"58",x"60",x"A9",x"00",x"8D",x"6C",x"02"
		,x"8D",x"6D",x"02",x"60",x"78",x"8A",x"48",x"A9"
		,x"50",x"8D",x"6C",x"02",x"A2",x"00",x"BD",x"CA"
		,x"FE",x"8D",x"6D",x"02",x"0D",x"00",x"1C",x"8D"
		,x"00",x"1C",x"68",x"AA",x"58",x"60",x"A9",x"00"
		,x"8D",x"F9",x"02",x"AD",x"8E",x"02",x"85",x"7F"
		,x"20",x"BC",x"E6",x"A5",x"84",x"10",x"09",x"29"
		,x"0F",x"C9",x"0F",x"F0",x"03",x"4C",x"B4",x"D7"
		,x"20",x"B3",x"C2",x"B1",x"A3",x"8D",x"75",x"02"
		,x"A2",x"0B",x"BD",x"89",x"FE",x"CD",x"75",x"02"
		,x"F0",x"08",x"CA",x"10",x"F5",x"A9",x"31",x"4C"
		,x"C8",x"C1",x"8E",x"2A",x"02",x"E0",x"09",x"90"
		,x"03",x"20",x"EE",x"C1",x"AE",x"2A",x"02",x"BD"
		,x"95",x"FE",x"85",x"6F",x"BD",x"A1",x"FE",x"85"
		,x"70",x"6C",x"6F",x"00",x"A9",x"00",x"8D",x"F9"
		,x"02",x"AD",x"6C",x"02",x"D0",x"2A",x"A0",x"00"
		,x"98",x"84",x"80",x"84",x"81",x"84",x"A3",x"20"
		,x"C7",x"E6",x"20",x"23",x"C1",x"A5",x"7F",x"8D"
		,x"8E",x"02",x"AA",x"4C",x"62",x"FF",x"EA",x"20"
		,x"BD",x"C1",x"4C",x"DA",x"D4",x"A0",x"28",x"A9"
		,x"00",x"99",x"00",x"02",x"88",x"10",x"FA",x"60"
		,x"A0",x"00",x"84",x"80",x"84",x"81",x"4C",x"45"
		,x"E6",x"A2",x"00",x"8E",x"7A",x"02",x"A9",x"3A"
		,x"20",x"68",x"C2",x"F0",x"05",x"88",x"88",x"8C"
		,x"7A",x"02",x"4C",x"68",x"C3",x"A0",x"00",x"A2"
		,x"00",x"A9",x"3A",x"4C",x"68",x"C2",x"20",x"E5"
		,x"C1",x"D0",x"05",x"A9",x"34",x"4C",x"C8",x"C1"
		,x"88",x"88",x"8C",x"7A",x"02",x"8A",x"D0",x"F3"
		,x"A9",x"3D",x"20",x"68",x"C2",x"8A",x"F0",x"02"
		,x"A9",x"40",x"09",x"21",x"8D",x"8B",x"02",x"E8"
		,x"8E",x"77",x"02",x"8E",x"78",x"02",x"AD",x"8A"
		,x"02",x"F0",x"0D",x"A9",x"80",x"0D",x"8B",x"02"
		,x"8D",x"8B",x"02",x"A9",x"00",x"8D",x"8A",x"02"
		,x"98",x"F0",x"29",x"9D",x"7A",x"02",x"AD",x"77"
		,x"02",x"8D",x"79",x"02",x"A9",x"8D",x"20",x"68"
		,x"C2",x"E8",x"8E",x"78",x"02",x"CA",x"AD",x"8A"
		,x"02",x"F0",x"02",x"A9",x"08",x"EC",x"77",x"02"
		,x"F0",x"02",x"09",x"04",x"09",x"03",x"4D",x"8B"
		,x"02",x"8D",x"8B",x"02",x"AD",x"8B",x"02",x"AE"
		,x"2A",x"02",x"3D",x"A5",x"FE",x"D0",x"01",x"60"
		,x"8D",x"6C",x"02",x"A9",x"30",x"4C",x"C8",x"C1"
		,x"8D",x"75",x"02",x"CC",x"74",x"02",x"B0",x"2E"
		,x"B1",x"A3",x"C8",x"CD",x"75",x"02",x"F0",x"28"
		,x"C9",x"2A",x"F0",x"04",x"C9",x"3F",x"D0",x"03"
		,x"EE",x"8A",x"02",x"C9",x"2C",x"D0",x"E4",x"98"
		,x"9D",x"7B",x"02",x"AD",x"8A",x"02",x"29",x"7F"
		,x"F0",x"07",x"A9",x"80",x"95",x"E7",x"8D",x"8A"
		,x"02",x"E8",x"E0",x"04",x"90",x"CD",x"A0",x"00"
		,x"AD",x"74",x"02",x"9D",x"7B",x"02",x"AD",x"8A"
		,x"02",x"29",x"7F",x"F0",x"04",x"A9",x"80",x"95"
		,x"E7",x"98",x"60",x"A4",x"A3",x"F0",x"14",x"88"
		,x"F0",x"10",x"B9",x"00",x"02",x"C9",x"0D",x"F0"
		,x"0A",x"88",x"B9",x"00",x"02",x"C9",x"0D",x"F0"
		,x"02",x"C8",x"C8",x"8C",x"74",x"02",x"C0",x"2A"
		,x"A0",x"FF",x"90",x"08",x"8C",x"2A",x"02",x"A9"
		,x"32",x"4C",x"C8",x"C1",x"A0",x"00",x"98",x"85"
		,x"A3",x"8D",x"58",x"02",x"8D",x"4A",x"02",x"8D"
		,x"96",x"02",x"85",x"D3",x"8D",x"79",x"02",x"8D"
		,x"77",x"02",x"8D",x"78",x"02",x"8D",x"8A",x"02"
		,x"8D",x"6C",x"02",x"A2",x"05",x"9D",x"79",x"02"
		,x"95",x"D7",x"95",x"DC",x"95",x"E1",x"95",x"E6"
		,x"9D",x"7F",x"02",x"9D",x"84",x"02",x"CA",x"D0"
		,x"EC",x"60",x"AD",x"78",x"02",x"8D",x"77",x"02"
		,x"A9",x"01",x"8D",x"78",x"02",x"8D",x"79",x"02"
		,x"AC",x"8E",x"02",x"A2",x"00",x"86",x"D3",x"BD"
		,x"7A",x"02",x"20",x"3C",x"C3",x"A6",x"D3",x"9D"
		,x"7A",x"02",x"98",x"95",x"E2",x"E8",x"EC",x"78"
		,x"02",x"90",x"EA",x"60",x"AA",x"A0",x"00",x"A9"
		,x"3A",x"DD",x"01",x"02",x"F0",x"0C",x"DD",x"00"
		,x"02",x"D0",x"16",x"E8",x"98",x"29",x"01",x"A8"
		,x"8A",x"60",x"BD",x"00",x"02",x"E8",x"E8",x"C9"
		,x"30",x"F0",x"F2",x"C9",x"31",x"F0",x"EE",x"D0"
		,x"EB",x"98",x"09",x"80",x"29",x"81",x"D0",x"E7"
		,x"A9",x"00",x"8D",x"8B",x"02",x"AC",x"7A",x"02"
		,x"B1",x"A3",x"20",x"BD",x"C3",x"10",x"11",x"C8"
		,x"CC",x"74",x"02",x"B0",x"06",x"AC",x"74",x"02"
		,x"88",x"D0",x"ED",x"CE",x"8B",x"02",x"A9",x"00"
		,x"29",x"01",x"85",x"7F",x"4C",x"00",x"C1",x"A5"
		,x"7F",x"49",x"01",x"29",x"01",x"85",x"7F",x"60"
		,x"A0",x"00",x"AD",x"77",x"02",x"CD",x"78",x"02"
		,x"F0",x"16",x"CE",x"78",x"02",x"AC",x"78",x"02"
		,x"B9",x"7A",x"02",x"A8",x"B1",x"A3",x"A0",x"04"
		,x"D9",x"BB",x"FE",x"F0",x"03",x"88",x"D0",x"F8"
		,x"98",x"8D",x"96",x"02",x"60",x"C9",x"30",x"F0"
		,x"06",x"C9",x"31",x"F0",x"02",x"09",x"80",x"29"
		,x"81",x"60",x"A9",x"00",x"85",x"6F",x"8D",x"8D"
		,x"02",x"48",x"AE",x"78",x"02",x"68",x"05",x"6F"
		,x"48",x"A9",x"01",x"85",x"6F",x"CA",x"30",x"0F"
		,x"B5",x"E2",x"10",x"04",x"06",x"6F",x"06",x"6F"
		,x"4A",x"90",x"EA",x"06",x"6F",x"D0",x"E6",x"68"
		,x"AA",x"BD",x"3F",x"C4",x"48",x"29",x"03",x"8D"
		,x"8C",x"02",x"68",x"0A",x"10",x"3E",x"A5",x"E2"
		,x"29",x"01",x"85",x"7F",x"AD",x"8C",x"02",x"F0"
		,x"2B",x"20",x"3D",x"C6",x"F0",x"12",x"20",x"8F"
		,x"C3",x"A9",x"00",x"8D",x"8C",x"02",x"20",x"3D"
		,x"C6",x"F0",x"1E",x"A9",x"74",x"20",x"C8",x"C1"
		,x"20",x"8F",x"C3",x"20",x"3D",x"C6",x"08",x"20"
		,x"8F",x"C3",x"28",x"F0",x"0C",x"A9",x"00",x"8D"
		,x"8C",x"02",x"F0",x"05",x"20",x"3D",x"C6",x"D0"
		,x"E2",x"4C",x"00",x"C1",x"2A",x"4C",x"00",x"C4"
		,x"00",x"80",x"41",x"01",x"01",x"01",x"01",x"81"
		,x"81",x"81",x"81",x"42",x"42",x"42",x"42",x"20"
		,x"CA",x"C3",x"A9",x"00",x"8D",x"92",x"02",x"20"
		,x"AC",x"C5",x"D0",x"19",x"CE",x"8C",x"02",x"10"
		,x"01",x"60",x"A9",x"01",x"8D",x"8D",x"02",x"20"
		,x"8F",x"C3",x"20",x"00",x"C1",x"4C",x"52",x"C4"
		,x"20",x"17",x"C6",x"F0",x"10",x"20",x"D8",x"C4"
		,x"AD",x"8F",x"02",x"F0",x"01",x"60",x"AD",x"53"
		,x"02",x"30",x"ED",x"10",x"F0",x"AD",x"8F",x"02"
		,x"F0",x"D2",x"60",x"20",x"04",x"C6",x"F0",x"1A"
		,x"D0",x"28",x"A9",x"01",x"8D",x"8D",x"02",x"20"
		,x"8F",x"C3",x"20",x"00",x"C1",x"A9",x"00",x"8D"
		,x"92",x"02",x"20",x"AC",x"C5",x"D0",x"13",x"8D"
		,x"8F",x"02",x"AD",x"8F",x"02",x"D0",x"28",x"CE"
		,x"8C",x"02",x"10",x"DE",x"60",x"20",x"17",x"C6"
		,x"F0",x"F0",x"20",x"D8",x"C4",x"AE",x"53",x"02"
		,x"10",x"07",x"AD",x"8F",x"02",x"F0",x"EE",x"D0"
		,x"0E",x"AD",x"96",x"02",x"F0",x"09",x"B5",x"E7"
		,x"29",x"07",x"CD",x"96",x"02",x"D0",x"DE",x"60"
		,x"A2",x"FF",x"8E",x"53",x"02",x"E8",x"8E",x"8A"
		,x"02",x"20",x"89",x"C5",x"F0",x"06",x"60",x"20"
		,x"94",x"C5",x"D0",x"FA",x"A5",x"7F",x"55",x"E2"
		,x"4A",x"90",x"0B",x"29",x"40",x"F0",x"F0",x"A9"
		,x"02",x"CD",x"8C",x"02",x"F0",x"E9",x"BD",x"7A"
		,x"02",x"AA",x"20",x"A6",x"C6",x"A0",x"03",x"4C"
		,x"1D",x"C5",x"BD",x"00",x"02",x"D1",x"94",x"F0"
		,x"0A",x"C9",x"3F",x"D0",x"D2",x"B1",x"94",x"C9"
		,x"A0",x"F0",x"CC",x"E8",x"C8",x"EC",x"76",x"02"
		,x"B0",x"09",x"BD",x"00",x"02",x"C9",x"2A",x"F0"
		,x"0C",x"D0",x"DF",x"C0",x"13",x"B0",x"06",x"B1"
		,x"94",x"C9",x"A0",x"D0",x"B2",x"AE",x"79",x"02"
		,x"8E",x"53",x"02",x"B5",x"E7",x"29",x"80",x"8D"
		,x"8A",x"02",x"AD",x"94",x"02",x"95",x"DD",x"A5"
		,x"81",x"95",x"D8",x"A0",x"00",x"B1",x"94",x"C8"
		,x"48",x"29",x"40",x"85",x"6F",x"68",x"29",x"DF"
		,x"30",x"02",x"09",x"20",x"29",x"27",x"05",x"6F"
		,x"85",x"6F",x"A9",x"80",x"35",x"E7",x"05",x"6F"
		,x"95",x"E7",x"B5",x"E2",x"29",x"80",x"05",x"7F"
		,x"95",x"E2",x"B1",x"94",x"9D",x"80",x"02",x"C8"
		,x"B1",x"94",x"9D",x"85",x"02",x"AD",x"58",x"02"
		,x"D0",x"07",x"A0",x"15",x"B1",x"94",x"8D",x"58"
		,x"02",x"A9",x"FF",x"8D",x"8F",x"02",x"AD",x"78"
		,x"02",x"8D",x"79",x"02",x"CE",x"79",x"02",x"10"
		,x"01",x"60",x"AE",x"79",x"02",x"B5",x"E7",x"30"
		,x"05",x"BD",x"80",x"02",x"D0",x"EE",x"A9",x"00"
		,x"8D",x"8F",x"02",x"60",x"A0",x"00",x"8C",x"91"
		,x"02",x"88",x"8C",x"53",x"02",x"AD",x"85",x"FE"
		,x"85",x"80",x"A9",x"01",x"85",x"81",x"8D",x"93"
		,x"02",x"20",x"75",x"D4",x"AD",x"93",x"02",x"D0"
		,x"01",x"60",x"A9",x"07",x"8D",x"95",x"02",x"A9"
		,x"00",x"20",x"F6",x"D4",x"8D",x"93",x"02",x"20"
		,x"E8",x"D4",x"CE",x"95",x"02",x"A0",x"00",x"B1"
		,x"94",x"D0",x"18",x"AD",x"91",x"02",x"D0",x"2F"
		,x"20",x"3B",x"DE",x"A5",x"81",x"8D",x"91",x"02"
		,x"A5",x"94",x"AE",x"92",x"02",x"8D",x"92",x"02"
		,x"F0",x"1D",x"60",x"A2",x"01",x"EC",x"92",x"02"
		,x"D0",x"2D",x"F0",x"13",x"AD",x"85",x"FE",x"85"
		,x"80",x"AD",x"90",x"02",x"85",x"81",x"20",x"75"
		,x"D4",x"AD",x"94",x"02",x"20",x"C8",x"D4",x"A9"
		,x"FF",x"8D",x"53",x"02",x"AD",x"95",x"02",x"30"
		,x"08",x"A9",x"20",x"20",x"C6",x"D1",x"4C",x"D7"
		,x"C5",x"20",x"4D",x"D4",x"4C",x"C4",x"C5",x"A5"
		,x"94",x"8D",x"94",x"02",x"20",x"3B",x"DE",x"A5"
		,x"81",x"8D",x"90",x"02",x"60",x"A5",x"68",x"D0"
		,x"28",x"A6",x"7F",x"56",x"1C",x"90",x"22",x"A9"
		,x"FF",x"8D",x"98",x"02",x"20",x"0E",x"D0",x"A0"
		,x"FF",x"C9",x"02",x"F0",x"0A",x"C9",x"03",x"F0"
		,x"06",x"C9",x"0F",x"F0",x"02",x"A0",x"00",x"A6"
		,x"7F",x"4C",x"6A",x"FF",x"D0",x"03",x"20",x"42"
		,x"D0",x"A6",x"7F",x"4C",x"56",x"FF",x"48",x"20"
		,x"A6",x"C6",x"20",x"88",x"C6",x"68",x"38",x"ED"
		,x"4B",x"02",x"AA",x"F0",x"0A",x"90",x"08",x"A9"
		,x"A0",x"91",x"94",x"C8",x"CA",x"D0",x"FA",x"60"
		,x"98",x"0A",x"A8",x"B9",x"99",x"00",x"85",x"94"
		,x"B9",x"9A",x"00",x"85",x"95",x"A0",x"00",x"BD"
		,x"00",x"02",x"91",x"94",x"C8",x"F0",x"06",x"E8"
		,x"EC",x"76",x"02",x"90",x"F2",x"60",x"A9",x"00"
		,x"8D",x"4B",x"02",x"8A",x"48",x"BD",x"00",x"02"
		,x"C9",x"2C",x"F0",x"14",x"C9",x"3D",x"F0",x"10"
		,x"EE",x"4B",x"02",x"E8",x"A9",x"0F",x"CD",x"4B"
		,x"02",x"90",x"05",x"EC",x"74",x"02",x"90",x"E5"
		,x"8E",x"76",x"02",x"68",x"AA",x"60",x"A5",x"83"
		,x"48",x"A5",x"82",x"48",x"20",x"DE",x"C6",x"68"
		,x"85",x"82",x"68",x"85",x"83",x"60",x"A9",x"11"
		,x"85",x"83",x"20",x"EB",x"D0",x"20",x"E8",x"D4"
		,x"AD",x"53",x"02",x"10",x"0A",x"AD",x"8D",x"02"
		,x"D0",x"0A",x"20",x"06",x"C8",x"18",x"60",x"AD"
		,x"8D",x"02",x"F0",x"1F",x"CE",x"8D",x"02",x"D0"
		,x"0D",x"CE",x"8D",x"02",x"20",x"8F",x"C3",x"20"
		,x"06",x"C8",x"38",x"4C",x"8F",x"C3",x"A9",x"00"
		,x"8D",x"73",x"02",x"8D",x"8D",x"02",x"20",x"B7"
		,x"C7",x"38",x"60",x"A2",x"18",x"A0",x"1D",x"B1"
		,x"94",x"8D",x"73",x"02",x"F0",x"02",x"A2",x"16"
		,x"88",x"B1",x"94",x"8D",x"72",x"02",x"E0",x"16"
		,x"F0",x"0A",x"C9",x"0A",x"90",x"06",x"CA",x"C9"
		,x"64",x"90",x"01",x"CA",x"20",x"AC",x"C7",x"B1"
		,x"94",x"48",x"0A",x"10",x"05",x"A9",x"3C",x"9D"
		,x"B2",x"02",x"68",x"29",x"0F",x"A8",x"B9",x"C5"
		,x"FE",x"9D",x"B1",x"02",x"CA",x"B9",x"C0",x"FE"
		,x"9D",x"B1",x"02",x"CA",x"B9",x"BB",x"FE",x"9D"
		,x"B1",x"02",x"CA",x"CA",x"B0",x"05",x"A9",x"2A"
		,x"9D",x"B2",x"02",x"A9",x"A0",x"9D",x"B1",x"02"
		,x"CA",x"A0",x"12",x"B1",x"94",x"9D",x"B1",x"02"
		,x"CA",x"88",x"C0",x"03",x"B0",x"F5",x"A9",x"22"
		,x"9D",x"B1",x"02",x"E8",x"E0",x"20",x"B0",x"0B"
		,x"BD",x"B1",x"02",x"C9",x"22",x"F0",x"04",x"C9"
		,x"A0",x"D0",x"F0",x"A9",x"22",x"9D",x"B1",x"02"
		,x"E8",x"E0",x"20",x"B0",x"0A",x"A9",x"7F",x"3D"
		,x"B1",x"02",x"9D",x"B1",x"02",x"10",x"F1",x"20"
		,x"B5",x"C4",x"38",x"60",x"A0",x"1B",x"A9",x"20"
		,x"99",x"B0",x"02",x"88",x"D0",x"FA",x"60",x"20"
		,x"19",x"F1",x"20",x"DF",x"F0",x"20",x"AC",x"C7"
		,x"A9",x"FF",x"85",x"6F",x"A6",x"7F",x"8E",x"72"
		,x"02",x"A9",x"00",x"8D",x"73",x"02",x"A6",x"F9"
		,x"BD",x"E0",x"FE",x"85",x"95",x"AD",x"88",x"FE"
		,x"85",x"94",x"A0",x"16",x"B1",x"94",x"C9",x"A0"
		,x"D0",x"0B",x"A9",x"31",x"2C",x"B1",x"94",x"C9"
		,x"A0",x"D0",x"02",x"A9",x"20",x"99",x"B3",x"02"
		,x"88",x"10",x"F2",x"A9",x"12",x"8D",x"B1",x"02"
		,x"A9",x"22",x"8D",x"B2",x"02",x"8D",x"C3",x"02"
		,x"A9",x"20",x"8D",x"C4",x"02",x"60",x"20",x"AC"
		,x"C7",x"A0",x"0B",x"B9",x"17",x"C8",x"99",x"B1"
		,x"02",x"88",x"10",x"F7",x"4C",x"4D",x"EF",x"42"
		,x"4C",x"4F",x"43",x"4B",x"53",x"20",x"46",x"52"
		,x"45",x"45",x"2E",x"20",x"98",x"C3",x"20",x"20"
		,x"C3",x"20",x"CA",x"C3",x"A9",x"00",x"85",x"86"
		,x"20",x"9D",x"C4",x"30",x"3D",x"20",x"B7",x"DD"
		,x"90",x"33",x"A0",x"00",x"B1",x"94",x"29",x"40"
		,x"D0",x"2B",x"20",x"B6",x"C8",x"A0",x"13",x"B1"
		,x"94",x"F0",x"0A",x"85",x"80",x"C8",x"B1",x"94"
		,x"85",x"81",x"20",x"7D",x"C8",x"AE",x"53",x"02"
		,x"A9",x"20",x"35",x"E7",x"D0",x"0D",x"BD",x"80"
		,x"02",x"85",x"80",x"BD",x"85",x"02",x"85",x"81"
		,x"20",x"7D",x"C8",x"E6",x"86",x"20",x"8B",x"C4"
		,x"10",x"C3",x"A5",x"86",x"85",x"80",x"A9",x"01"
		,x"A0",x"00",x"4C",x"A3",x"C1",x"20",x"5F",x"EF"
		,x"20",x"75",x"D4",x"20",x"19",x"F1",x"B5",x"A7"
		,x"C9",x"FF",x"F0",x"08",x"AD",x"F9",x"02",x"09"
		,x"40",x"8D",x"F9",x"02",x"A9",x"00",x"20",x"C8"
		,x"D4",x"20",x"56",x"D1",x"85",x"80",x"20",x"56"
		,x"D1",x"85",x"81",x"A5",x"80",x"D0",x"06",x"20"
		,x"F4",x"EE",x"4C",x"27",x"D2",x"20",x"5F",x"EF"
		,x"20",x"4D",x"D4",x"4C",x"94",x"C8",x"A0",x"00"
		,x"98",x"91",x"94",x"20",x"5E",x"DE",x"4C",x"99"
		,x"D5",x"A9",x"31",x"4C",x"C8",x"C1",x"A9",x"4C"
		,x"8D",x"00",x"06",x"A9",x"C7",x"8D",x"01",x"06"
		,x"A9",x"FA",x"8D",x"02",x"06",x"A9",x"03",x"20"
		,x"D3",x"D6",x"A5",x"7F",x"09",x"E0",x"85",x"03"
		,x"A5",x"03",x"30",x"FC",x"C9",x"02",x"90",x"07"
		,x"A9",x"03",x"A2",x"00",x"4C",x"0A",x"E6",x"60"
		,x"A9",x"E0",x"8D",x"4F",x"02",x"20",x"D1",x"F0"
		,x"20",x"19",x"F1",x"A9",x"FF",x"95",x"A7",x"A9"
		,x"0F",x"8D",x"56",x"02",x"20",x"E5",x"C1",x"D0"
		,x"03",x"4C",x"C1",x"C8",x"20",x"F8",x"C1",x"20"
		,x"20",x"C3",x"AD",x"8B",x"02",x"29",x"55",x"D0"
		,x"0F",x"AE",x"7A",x"02",x"BD",x"00",x"02",x"C9"
		,x"2A",x"D0",x"05",x"A9",x"30",x"4C",x"C8",x"C1"
		,x"AD",x"8B",x"02",x"29",x"D9",x"D0",x"F4",x"4C"
		,x"52",x"C9",x"A9",x"00",x"8D",x"58",x"02",x"8D"
		,x"8C",x"02",x"8D",x"80",x"02",x"8D",x"81",x"02"
		,x"A5",x"E3",x"29",x"01",x"85",x"7F",x"09",x"01"
		,x"8D",x"91",x"02",x"AD",x"7B",x"02",x"8D",x"7A"
		,x"02",x"60",x"20",x"4F",x"C4",x"AD",x"78",x"02"
		,x"C9",x"03",x"90",x"45",x"A5",x"E2",x"C5",x"E3"
		,x"D0",x"3F",x"A5",x"DD",x"C5",x"DE",x"D0",x"39"
		,x"A5",x"D8",x"C5",x"D9",x"D0",x"33",x"20",x"CC"
		,x"CA",x"A9",x"01",x"8D",x"79",x"02",x"20",x"FA"
		,x"C9",x"20",x"25",x"D1",x"F0",x"04",x"C9",x"02"
		,x"D0",x"05",x"A9",x"64",x"20",x"C8",x"C1",x"A9"
		,x"12",x"85",x"83",x"AD",x"3C",x"02",x"8D",x"3D"
		,x"02",x"A9",x"FF",x"8D",x"3C",x"02",x"20",x"2A"
		,x"DA",x"A2",x"02",x"20",x"B9",x"C9",x"4C",x"94"
		,x"C1",x"20",x"A7",x"C9",x"4C",x"94",x"C1",x"20"
		,x"E7",x"CA",x"A5",x"E2",x"29",x"01",x"85",x"7F"
		,x"20",x"86",x"D4",x"20",x"E4",x"D6",x"AE",x"77"
		,x"02",x"8E",x"79",x"02",x"20",x"FA",x"C9",x"A9"
		,x"11",x"85",x"83",x"20",x"EB",x"D0",x"20",x"25"
		,x"D1",x"D0",x"03",x"20",x"53",x"CA",x"A9",x"08"
		,x"85",x"F8",x"4C",x"D8",x"C9",x"20",x"9B",x"CF"
		,x"20",x"35",x"CA",x"A9",x"80",x"20",x"A6",x"DD"
		,x"F0",x"F3",x"20",x"25",x"D1",x"F0",x"03",x"20"
		,x"9B",x"CF",x"AE",x"79",x"02",x"E8",x"EC",x"78"
		,x"02",x"90",x"C6",x"A9",x"12",x"85",x"83",x"4C"
		,x"02",x"DB",x"AE",x"79",x"02",x"B5",x"E2",x"29"
		,x"01",x"85",x"7F",x"AD",x"85",x"FE",x"85",x"80"
		,x"B5",x"D8",x"85",x"81",x"20",x"75",x"D4",x"AE"
		,x"79",x"02",x"B5",x"DD",x"20",x"C8",x"D4",x"AE"
		,x"79",x"02",x"B5",x"E7",x"29",x"07",x"8D",x"4A"
		,x"02",x"A9",x"00",x"8D",x"58",x"02",x"20",x"A0"
		,x"D9",x"A0",x"01",x"20",x"25",x"D1",x"F0",x"01"
		,x"C8",x"98",x"4C",x"C8",x"D4",x"A9",x"11",x"85"
		,x"83",x"20",x"9B",x"D3",x"85",x"85",x"A6",x"82"
		,x"B5",x"F2",x"29",x"08",x"85",x"F8",x"D0",x"0A"
		,x"20",x"25",x"D1",x"F0",x"05",x"A9",x"80",x"20"
		,x"97",x"DD",x"60",x"20",x"D3",x"D1",x"20",x"CB"
		,x"E1",x"A5",x"D6",x"48",x"A5",x"D5",x"48",x"A9"
		,x"12",x"85",x"83",x"20",x"07",x"D1",x"20",x"D3"
		,x"D1",x"20",x"CB",x"E1",x"20",x"9C",x"E2",x"A5"
		,x"D6",x"85",x"87",x"A5",x"D5",x"85",x"86",x"A9"
		,x"00",x"85",x"88",x"85",x"D4",x"85",x"D7",x"68"
		,x"85",x"D5",x"68",x"85",x"D6",x"4C",x"3B",x"E3"
		,x"20",x"20",x"C3",x"A5",x"E3",x"29",x"01",x"85"
		,x"E3",x"C5",x"E2",x"F0",x"02",x"09",x"80",x"85"
		,x"E2",x"20",x"4F",x"C4",x"20",x"E7",x"CA",x"A5"
		,x"E3",x"29",x"01",x"85",x"7F",x"A5",x"D9",x"85"
		,x"81",x"20",x"57",x"DE",x"20",x"99",x"D5",x"A5"
		,x"DE",x"18",x"69",x"03",x"20",x"C8",x"D4",x"20"
		,x"93",x"DF",x"A8",x"AE",x"7A",x"02",x"A9",x"10"
		,x"20",x"6E",x"C6",x"20",x"5E",x"DE",x"20",x"99"
		,x"D5",x"4C",x"94",x"C1",x"A5",x"E8",x"29",x"07"
		,x"8D",x"4A",x"02",x"AE",x"78",x"02",x"CA",x"EC"
		,x"77",x"02",x"90",x"0A",x"BD",x"80",x"02",x"D0"
		,x"F5",x"A9",x"62",x"4C",x"C8",x"C1",x"60",x"20"
		,x"CC",x"CA",x"BD",x"80",x"02",x"F0",x"05",x"A9"
		,x"63",x"4C",x"C8",x"C1",x"CA",x"10",x"F3",x"60"
		,x"AD",x"01",x"02",x"C9",x"2D",x"D0",x"4C",x"AD"
		,x"03",x"02",x"85",x"6F",x"AD",x"04",x"02",x"85"
		,x"70",x"A0",x"00",x"AD",x"02",x"02",x"C9",x"52"
		,x"F0",x"0E",x"20",x"58",x"F2",x"C9",x"57",x"F0"
		,x"37",x"C9",x"45",x"D0",x"2E",x"6C",x"6F",x"00"
		,x"B1",x"6F",x"85",x"85",x"AD",x"74",x"02",x"C9"
		,x"06",x"90",x"1A",x"AE",x"05",x"02",x"CA",x"F0"
		,x"14",x"8A",x"18",x"65",x"6F",x"E6",x"6F",x"8D"
		,x"49",x"02",x"A5",x"6F",x"85",x"A5",x"A5",x"70"
		,x"85",x"A6",x"4C",x"43",x"D4",x"20",x"EB",x"D0"
		,x"4C",x"3A",x"D4",x"A9",x"31",x"4C",x"C8",x"C1"
		,x"B9",x"06",x"02",x"91",x"6F",x"C8",x"CC",x"05"
		,x"02",x"90",x"F5",x"60",x"AC",x"01",x"02",x"C0"
		,x"30",x"D0",x"09",x"A9",x"EA",x"85",x"6B",x"A9"
		,x"FF",x"85",x"6C",x"60",x"20",x"72",x"CB",x"4C"
		,x"94",x"C1",x"88",x"98",x"29",x"0F",x"0A",x"A8"
		,x"B1",x"6B",x"85",x"75",x"C8",x"B1",x"6B",x"85"
		,x"76",x"6C",x"75",x"00",x"AD",x"8E",x"02",x"85"
		,x"7F",x"A5",x"83",x"48",x"20",x"3D",x"C6",x"68"
		,x"85",x"83",x"AE",x"74",x"02",x"CA",x"D0",x"0D"
		,x"A9",x"01",x"20",x"E2",x"D1",x"4C",x"F1",x"CB"
		,x"A9",x"70",x"4C",x"C8",x"C1",x"A0",x"01",x"20"
		,x"7C",x"CC",x"AE",x"85",x"02",x"E0",x"05",x"B0"
		,x"EF",x"A9",x"00",x"85",x"6F",x"85",x"70",x"38"
		,x"26",x"6F",x"26",x"70",x"CA",x"10",x"F9",x"A5"
		,x"6F",x"2D",x"4F",x"02",x"D0",x"DA",x"A5",x"70"
		,x"2D",x"50",x"02",x"D0",x"D3",x"A5",x"6F",x"0D"
		,x"4F",x"02",x"8D",x"4F",x"02",x"A5",x"70",x"0D"
		,x"50",x"02",x"8D",x"50",x"02",x"A9",x"00",x"20"
		,x"E2",x"D1",x"A6",x"82",x"AD",x"85",x"02",x"95"
		,x"A7",x"AA",x"A5",x"7F",x"95",x"00",x"9D",x"5B"
		,x"02",x"A6",x"83",x"BD",x"2B",x"02",x"09",x"40"
		,x"9D",x"2B",x"02",x"A4",x"82",x"A9",x"FF",x"99"
		,x"44",x"02",x"A9",x"89",x"99",x"F2",x"00",x"B9"
		,x"A7",x"00",x"99",x"3E",x"02",x"0A",x"AA",x"A9"
		,x"01",x"95",x"99",x"A9",x"0E",x"99",x"EC",x"00"
		,x"4C",x"94",x"C1",x"A0",x"00",x"A2",x"00",x"A9"
		,x"2D",x"20",x"68",x"C2",x"D0",x"0A",x"A9",x"31"
		,x"4C",x"C8",x"C1",x"A9",x"30",x"4C",x"C8",x"C1"
		,x"8A",x"D0",x"F8",x"A2",x"05",x"B9",x"00",x"02"
		,x"DD",x"5D",x"CC",x"F0",x"05",x"CA",x"10",x"F8"
		,x"30",x"E4",x"8A",x"09",x"80",x"8D",x"2A",x"02"
		,x"20",x"6F",x"CC",x"AD",x"2A",x"02",x"0A",x"AA"
		,x"BD",x"64",x"CC",x"85",x"70",x"BD",x"63",x"CC"
		,x"85",x"6F",x"6C",x"6F",x"00",x"41",x"46",x"52"
		,x"57",x"45",x"50",x"03",x"CD",x"F5",x"CC",x"56"
		,x"CD",x"73",x"CD",x"A3",x"CD",x"BD",x"CD",x"A0"
		,x"00",x"A2",x"00",x"A9",x"3A",x"20",x"68",x"C2"
		,x"D0",x"02",x"A0",x"03",x"B9",x"00",x"02",x"C9"
		,x"20",x"F0",x"08",x"C9",x"1D",x"F0",x"04",x"C9"
		,x"2C",x"D0",x"07",x"C8",x"CC",x"74",x"02",x"90"
		,x"EB",x"60",x"20",x"A1",x"CC",x"EE",x"77",x"02"
		,x"AC",x"79",x"02",x"E0",x"04",x"90",x"EC",x"B0"
		,x"8A",x"A9",x"00",x"85",x"6F",x"85",x"70",x"85"
		,x"72",x"A2",x"FF",x"B9",x"00",x"02",x"C9",x"40"
		,x"B0",x"18",x"C9",x"30",x"90",x"14",x"29",x"0F"
		,x"48",x"A5",x"70",x"85",x"71",x"A5",x"6F",x"85"
		,x"70",x"68",x"85",x"6F",x"C8",x"CC",x"74",x"02"
		,x"90",x"E1",x"8C",x"79",x"02",x"18",x"A9",x"00"
		,x"E8",x"E0",x"03",x"B0",x"0F",x"B4",x"6F",x"88"
		,x"30",x"F6",x"7D",x"F2",x"CC",x"90",x"F8",x"18"
		,x"E6",x"72",x"D0",x"F3",x"48",x"AE",x"77",x"02"
		,x"A5",x"72",x"9D",x"80",x"02",x"68",x"9D",x"85"
		,x"02",x"60",x"01",x"0A",x"64",x"20",x"F5",x"CD"
		,x"20",x"5F",x"EF",x"4C",x"94",x"C1",x"A9",x"01"
		,x"8D",x"F9",x"02",x"20",x"F5",x"CD",x"A5",x"81"
		,x"48",x"20",x"FA",x"F1",x"F0",x"0B",x"68",x"C5"
		,x"81",x"D0",x"19",x"20",x"90",x"EF",x"4C",x"94"
		,x"C1",x"68",x"A9",x"00",x"85",x"81",x"E6",x"80"
		,x"A5",x"80",x"CD",x"D7",x"FE",x"B0",x"0A",x"20"
		,x"FA",x"F1",x"F0",x"EE",x"A9",x"65",x"20",x"45"
		,x"E6",x"A9",x"65",x"20",x"C8",x"C1",x"20",x"F2"
		,x"CD",x"4C",x"60",x"D4",x"20",x"2F",x"D1",x"A1"
		,x"99",x"60",x"20",x"36",x"CD",x"A9",x"00",x"20"
		,x"C8",x"D4",x"20",x"3C",x"CD",x"99",x"44",x"02"
		,x"A9",x"89",x"99",x"F2",x"00",x"60",x"20",x"42"
		,x"CD",x"20",x"EC",x"D3",x"4C",x"94",x"C1",x"20"
		,x"6F",x"CC",x"20",x"42",x"CD",x"B9",x"44",x"02"
		,x"99",x"3E",x"02",x"A9",x"FF",x"99",x"44",x"02"
		,x"4C",x"94",x"C1",x"20",x"F2",x"CD",x"20",x"E8"
		,x"D4",x"A8",x"88",x"C9",x"02",x"B0",x"02",x"A0"
		,x"01",x"A9",x"00",x"20",x"C8",x"D4",x"98",x"20"
		,x"F1",x"CF",x"8A",x"48",x"20",x"64",x"D4",x"68"
		,x"AA",x"20",x"70",x"C0",x"4C",x"94",x"C1",x"20"
		,x"6F",x"CC",x"20",x"F2",x"CD",x"20",x"64",x"D4"
		,x"4C",x"94",x"C1",x"20",x"58",x"F2",x"20",x"36"
		,x"CD",x"A9",x"00",x"85",x"6F",x"A6",x"F9",x"BD"
		,x"E0",x"FE",x"85",x"70",x"20",x"BA",x"CD",x"4C"
		,x"94",x"C1",x"6C",x"6F",x"00",x"20",x"D2",x"CD"
		,x"A5",x"F9",x"0A",x"AA",x"AD",x"86",x"02",x"95"
		,x"99",x"20",x"2F",x"D1",x"20",x"EE",x"D3",x"4C"
		,x"94",x"C1",x"A6",x"D3",x"E6",x"D3",x"BD",x"85"
		,x"02",x"A8",x"88",x"88",x"C0",x"0C",x"90",x"05"
		,x"A9",x"70",x"4C",x"C8",x"C1",x"85",x"83",x"20"
		,x"EB",x"D0",x"B0",x"F4",x"20",x"93",x"DF",x"85"
		,x"F9",x"60",x"20",x"D2",x"CD",x"A6",x"D3",x"BD"
		,x"85",x"02",x"29",x"01",x"85",x"7F",x"BD",x"87"
		,x"02",x"85",x"81",x"BD",x"86",x"02",x"85",x"80"
		,x"20",x"5F",x"D5",x"4C",x"00",x"C1",x"20",x"2C"
		,x"CE",x"20",x"6E",x"CE",x"A5",x"90",x"85",x"D7"
		,x"20",x"71",x"CE",x"E6",x"D7",x"E6",x"D7",x"A5"
		,x"8B",x"85",x"D5",x"A5",x"90",x"0A",x"18",x"69"
		,x"10",x"85",x"D6",x"60",x"20",x"D9",x"CE",x"85"
		,x"92",x"A6",x"82",x"B5",x"B5",x"85",x"90",x"B5"
		,x"BB",x"85",x"91",x"D0",x"04",x"A5",x"90",x"F0"
		,x"0B",x"A5",x"90",x"38",x"E9",x"01",x"85",x"90"
		,x"B0",x"02",x"C6",x"91",x"B5",x"C7",x"85",x"6F"
		,x"46",x"6F",x"90",x"03",x"20",x"ED",x"CE",x"20"
		,x"E5",x"CE",x"A5",x"6F",x"D0",x"F2",x"A5",x"D4"
		,x"18",x"65",x"8B",x"85",x"8B",x"90",x"06",x"E6"
		,x"8C",x"D0",x"02",x"E6",x"8D",x"60",x"A9",x"FE"
		,x"2C",x"A9",x"78",x"85",x"6F",x"A2",x"03",x"B5"
		,x"8F",x"48",x"B5",x"8A",x"95",x"8F",x"68",x"95"
		,x"8A",x"CA",x"D0",x"F3",x"20",x"D9",x"CE",x"A2"
		,x"00",x"B5",x"90",x"95",x"8F",x"E8",x"E0",x"04"
		,x"90",x"F7",x"A9",x"00",x"85",x"92",x"24",x"6F"
		,x"30",x"09",x"06",x"8F",x"08",x"46",x"8F",x"28"
		,x"20",x"E6",x"CE",x"20",x"ED",x"CE",x"20",x"E5"
		,x"CE",x"24",x"6F",x"30",x"03",x"20",x"E2",x"CE"
		,x"A5",x"8F",x"18",x"65",x"90",x"85",x"90",x"90"
		,x"06",x"E6",x"91",x"D0",x"02",x"E6",x"92",x"A5"
		,x"92",x"05",x"91",x"D0",x"C2",x"A5",x"90",x"38"
		,x"E5",x"6F",x"90",x"0C",x"E6",x"8B",x"D0",x"06"
		,x"E6",x"8C",x"D0",x"02",x"E6",x"8D",x"85",x"90"
		,x"60",x"A9",x"00",x"85",x"8B",x"85",x"8C",x"85"
		,x"8D",x"60",x"20",x"E5",x"CE",x"18",x"26",x"90"
		,x"26",x"91",x"26",x"92",x"60",x"18",x"A2",x"FD"
		,x"B5",x"8E",x"75",x"93",x"95",x"8E",x"E8",x"D0"
		,x"F7",x"60",x"A2",x"00",x"8A",x"95",x"FA",x"E8"
		,x"E0",x"04",x"D0",x"F8",x"A9",x"06",x"95",x"FA"
		,x"60",x"A0",x"04",x"A6",x"82",x"B9",x"FA",x"00"
		,x"96",x"FA",x"C5",x"82",x"F0",x"07",x"88",x"30"
		,x"E1",x"AA",x"4C",x"0D",x"CF",x"60",x"20",x"09"
		,x"CF",x"20",x"B7",x"DF",x"D0",x"46",x"20",x"D3"
		,x"D1",x"20",x"8E",x"D2",x"30",x"48",x"20",x"C2"
		,x"DF",x"A5",x"80",x"48",x"A5",x"81",x"48",x"A9"
		,x"01",x"20",x"F6",x"D4",x"85",x"81",x"A9",x"00"
		,x"20",x"F6",x"D4",x"85",x"80",x"F0",x"1F",x"20"
		,x"25",x"D1",x"F0",x"0B",x"20",x"AB",x"DD",x"D0"
		,x"06",x"20",x"8C",x"CF",x"4C",x"5D",x"CF",x"20"
		,x"8C",x"CF",x"20",x"57",x"DE",x"68",x"85",x"81"
		,x"68",x"85",x"80",x"4C",x"6F",x"CF",x"68",x"85"
		,x"81",x"68",x"85",x"80",x"20",x"8C",x"CF",x"20"
		,x"93",x"DF",x"AA",x"4C",x"99",x"D5",x"A9",x"70"
		,x"4C",x"C8",x"C1",x"20",x"09",x"CF",x"20",x"B7"
		,x"DF",x"D0",x"08",x"20",x"8E",x"D2",x"30",x"EE"
		,x"20",x"C2",x"DF",x"60",x"A6",x"82",x"B5",x"A7"
		,x"49",x"80",x"95",x"A7",x"B5",x"AE",x"49",x"80"
		,x"95",x"AE",x"60",x"A2",x"12",x"86",x"83",x"20"
		,x"07",x"D1",x"20",x"00",x"C1",x"20",x"25",x"D1"
		,x"90",x"05",x"A9",x"20",x"20",x"9D",x"DD",x"A5"
		,x"83",x"C9",x"0F",x"F0",x"23",x"D0",x"08",x"A5"
		,x"84",x"29",x"8F",x"C9",x"0F",x"B0",x"19",x"20"
		,x"25",x"D1",x"B0",x"05",x"A5",x"85",x"4C",x"9D"
		,x"D1",x"D0",x"03",x"4C",x"AB",x"E0",x"A5",x"85"
		,x"20",x"F1",x"CF",x"A4",x"82",x"4C",x"EE",x"D3"
		,x"A9",x"04",x"85",x"82",x"20",x"E8",x"D4",x"C9"
		,x"2A",x"F0",x"05",x"A5",x"85",x"20",x"F1",x"CF"
		,x"A5",x"F8",x"F0",x"01",x"60",x"EE",x"55",x"02"
		,x"60",x"48",x"20",x"93",x"DF",x"10",x"06",x"68"
		,x"A9",x"61",x"4C",x"C8",x"C1",x"0A",x"AA",x"68"
		,x"81",x"99",x"F6",x"99",x"60",x"20",x"D1",x"C1"
		,x"20",x"42",x"D0",x"4C",x"94",x"C1",x"20",x"0F"
		,x"F1",x"A8",x"B6",x"A7",x"E0",x"FF",x"D0",x"14"
		,x"48",x"20",x"8E",x"D2",x"AA",x"10",x"05",x"A9"
		,x"70",x"20",x"48",x"E6",x"68",x"A8",x"8A",x"09"
		,x"80",x"99",x"A7",x"00",x"8A",x"29",x"0F",x"85"
		,x"F9",x"A2",x"00",x"86",x"81",x"AE",x"85",x"FE"
		,x"86",x"80",x"20",x"D3",x"D6",x"A9",x"B0",x"4C"
		,x"8C",x"D5",x"20",x"D1",x"F0",x"20",x"13",x"D3"
		,x"20",x"0E",x"D0",x"A6",x"7F",x"A9",x"00",x"9D"
		,x"51",x"02",x"8A",x"0A",x"AA",x"A5",x"16",x"95"
		,x"12",x"A5",x"17",x"95",x"13",x"20",x"86",x"D5"
		,x"A5",x"F9",x"0A",x"AA",x"A9",x"02",x"95",x"99"
		,x"A1",x"99",x"A6",x"7F",x"9D",x"01",x"01",x"A9"
		,x"00",x"4C",x"71",x"FF",x"EA",x"20",x"3A",x"EF"
		,x"A0",x"04",x"A9",x"00",x"AA",x"18",x"71",x"6D"
		,x"90",x"01",x"E8",x"C8",x"C8",x"C8",x"C8",x"C0"
		,x"48",x"F0",x"F8",x"C0",x"90",x"D0",x"EE",x"48"
		,x"8A",x"A6",x"7F",x"9D",x"FC",x"02",x"68",x"9D"
		,x"FA",x"02",x"60",x"20",x"D0",x"D6",x"20",x"C3"
		,x"D0",x"20",x"99",x"D5",x"20",x"37",x"D1",x"85"
		,x"80",x"20",x"37",x"D1",x"85",x"81",x"60",x"20"
		,x"9B",x"D0",x"A5",x"80",x"D0",x"01",x"60",x"20"
		,x"1E",x"CF",x"20",x"D0",x"D6",x"20",x"C3",x"D0"
		,x"4C",x"1E",x"CF",x"A9",x"80",x"D0",x"02",x"A9"
		,x"90",x"8D",x"4D",x"02",x"20",x"93",x"DF",x"AA"
		,x"20",x"06",x"D5",x"8A",x"48",x"0A",x"AA",x"A9"
		,x"00",x"95",x"99",x"20",x"25",x"D1",x"C9",x"04"
		,x"B0",x"06",x"F6",x"B5",x"D0",x"02",x"F6",x"BB"
		,x"68",x"AA",x"60",x"A5",x"83",x"C9",x"13",x"90"
		,x"02",x"29",x"0F",x"C9",x"0F",x"D0",x"02",x"A9"
		,x"10",x"AA",x"38",x"BD",x"2B",x"02",x"30",x"06"
		,x"29",x"0F",x"85",x"82",x"AA",x"18",x"60",x"A5"
		,x"83",x"C9",x"13",x"90",x"02",x"29",x"0F",x"AA"
		,x"BD",x"2B",x"02",x"A8",x"0A",x"90",x"0A",x"30"
		,x"0A",x"98",x"29",x"0F",x"85",x"82",x"AA",x"18"
		,x"60",x"30",x"F6",x"38",x"60",x"A6",x"82",x"B5"
		,x"EC",x"4A",x"29",x"07",x"C9",x"04",x"60",x"20"
		,x"93",x"DF",x"0A",x"AA",x"A4",x"82",x"60",x"20"
		,x"2F",x"D1",x"B9",x"44",x"02",x"F0",x"12",x"A1"
		,x"99",x"48",x"B5",x"99",x"D9",x"44",x"02",x"D0"
		,x"04",x"A9",x"FF",x"95",x"99",x"68",x"F6",x"99"
		,x"60",x"A1",x"99",x"F6",x"99",x"60",x"20",x"37"
		,x"D1",x"D0",x"36",x"85",x"85",x"B9",x"44",x"02"
		,x"F0",x"08",x"A9",x"80",x"99",x"F2",x"00",x"A5"
		,x"85",x"60",x"20",x"1E",x"CF",x"A9",x"00",x"20"
		,x"C8",x"D4",x"20",x"37",x"D1",x"C9",x"00",x"F0"
		,x"19",x"85",x"80",x"20",x"37",x"D1",x"85",x"81"
		,x"20",x"1E",x"CF",x"20",x"D3",x"D1",x"20",x"D0"
		,x"D6",x"20",x"C3",x"D0",x"20",x"1E",x"CF",x"A5"
		,x"85",x"60",x"20",x"37",x"D1",x"A4",x"82",x"99"
		,x"44",x"02",x"A5",x"85",x"60",x"20",x"F1",x"CF"
		,x"F0",x"01",x"60",x"20",x"D3",x"D1",x"20",x"1E"
		,x"F1",x"A9",x"00",x"20",x"C8",x"D4",x"A5",x"80"
		,x"20",x"F1",x"CF",x"A5",x"81",x"20",x"F1",x"CF"
		,x"20",x"C7",x"D0",x"20",x"1E",x"CF",x"20",x"D0"
		,x"D6",x"A9",x"02",x"4C",x"C8",x"D4",x"85",x"6F"
		,x"20",x"E8",x"D4",x"18",x"65",x"6F",x"95",x"99"
		,x"85",x"94",x"60",x"20",x"93",x"DF",x"AA",x"BD"
		,x"5B",x"02",x"29",x"01",x"85",x"7F",x"60",x"38"
		,x"B0",x"01",x"18",x"08",x"85",x"6F",x"20",x"27"
		,x"D2",x"20",x"7F",x"D3",x"85",x"82",x"A6",x"83"
		,x"28",x"90",x"02",x"09",x"80",x"9D",x"2B",x"02"
		,x"29",x"3F",x"A8",x"A9",x"FF",x"99",x"A7",x"00"
		,x"99",x"AE",x"00",x"99",x"CD",x"00",x"C6",x"6F"
		,x"30",x"1C",x"20",x"8E",x"D2",x"10",x"08",x"20"
		,x"5A",x"D2",x"A9",x"70",x"4C",x"C8",x"C1",x"99"
		,x"A7",x"00",x"C6",x"6F",x"30",x"08",x"20",x"8E"
		,x"D2",x"30",x"EC",x"99",x"AE",x"00",x"60",x"A5"
		,x"83",x"C9",x"0F",x"D0",x"01",x"60",x"A6",x"83"
		,x"BD",x"2B",x"02",x"C9",x"FF",x"F0",x"22",x"29"
		,x"3F",x"85",x"82",x"A9",x"FF",x"9D",x"2B",x"02"
		,x"A6",x"82",x"A9",x"00",x"95",x"F2",x"20",x"5A"
		,x"D2",x"A6",x"82",x"A9",x"01",x"CA",x"30",x"03"
		,x"0A",x"D0",x"FA",x"0D",x"56",x"02",x"8D",x"56"
		,x"02",x"60",x"A6",x"82",x"B5",x"A7",x"C9",x"FF"
		,x"F0",x"09",x"48",x"A9",x"FF",x"95",x"A7",x"68"
		,x"20",x"F3",x"D2",x"A6",x"82",x"B5",x"AE",x"C9"
		,x"FF",x"F0",x"09",x"48",x"A9",x"FF",x"95",x"AE"
		,x"68",x"20",x"F3",x"D2",x"A6",x"82",x"B5",x"CD"
		,x"C9",x"FF",x"F0",x"09",x"48",x"A9",x"FF",x"95"
		,x"CD",x"68",x"20",x"F3",x"D2",x"60",x"98",x"48"
		,x"A0",x"01",x"20",x"BA",x"D2",x"10",x"0C",x"88"
		,x"20",x"BA",x"D2",x"10",x"06",x"20",x"39",x"D3"
		,x"AA",x"30",x"13",x"B5",x"00",x"30",x"FC",x"A5"
		,x"7F",x"95",x"00",x"9D",x"5B",x"02",x"8A",x"0A"
		,x"A8",x"A9",x"02",x"99",x"99",x"00",x"68",x"A8"
		,x"8A",x"60",x"A2",x"07",x"B9",x"4F",x"02",x"3D"
		,x"E9",x"EF",x"F0",x"04",x"CA",x"10",x"F5",x"60"
		,x"B9",x"4F",x"02",x"5D",x"E9",x"EF",x"99",x"4F"
		,x"02",x"8A",x"88",x"30",x"03",x"18",x"69",x"08"
		,x"AA",x"60",x"A6",x"82",x"B5",x"A7",x"30",x"09"
		,x"8A",x"18",x"69",x"07",x"AA",x"B5",x"A7",x"10"
		,x"F0",x"C9",x"FF",x"F0",x"EC",x"48",x"A9",x"FF"
		,x"95",x"A7",x"68",x"29",x"0F",x"A8",x"C8",x"A2"
		,x"10",x"6E",x"50",x"02",x"6E",x"4F",x"02",x"88"
		,x"D0",x"01",x"18",x"CA",x"10",x"F3",x"60",x"A9"
		,x"0E",x"85",x"83",x"20",x"27",x"D2",x"C6",x"83"
		,x"D0",x"F9",x"60",x"A9",x"0E",x"85",x"83",x"A6"
		,x"83",x"BD",x"2B",x"02",x"C9",x"FF",x"F0",x"14"
		,x"29",x"3F",x"85",x"82",x"20",x"93",x"DF",x"AA"
		,x"BD",x"5B",x"02",x"29",x"01",x"C5",x"7F",x"D0"
		,x"03",x"20",x"27",x"D2",x"C6",x"83",x"10",x"DF"
		,x"60",x"A5",x"6F",x"48",x"A0",x"00",x"B6",x"FA"
		,x"B5",x"A7",x"10",x"04",x"C9",x"FF",x"D0",x"16"
		,x"8A",x"18",x"69",x"07",x"AA",x"B5",x"A7",x"10"
		,x"04",x"C9",x"FF",x"D0",x"09",x"C8",x"C0",x"05"
		,x"90",x"E4",x"A2",x"FF",x"D0",x"1C",x"86",x"6F"
		,x"29",x"3F",x"AA",x"B5",x"00",x"30",x"FC",x"4C"
		,x"3B",x"FF",x"EA",x"A6",x"6F",x"E0",x"07",x"90"
		,x"D7",x"B0",x"E2",x"A4",x"6F",x"A9",x"FF",x"99"
		,x"A7",x"00",x"68",x"85",x"6F",x"8A",x"60",x"A0"
		,x"00",x"A9",x"01",x"2C",x"56",x"02",x"D0",x"09"
		,x"C8",x"0A",x"D0",x"F7",x"A9",x"70",x"4C",x"C8"
		,x"C1",x"49",x"FF",x"2D",x"56",x"02",x"8D",x"56"
		,x"02",x"98",x"60",x"20",x"EB",x"D0",x"20",x"00"
		,x"C1",x"20",x"AA",x"D3",x"A6",x"82",x"BD",x"3E"
		,x"02",x"60",x"A6",x"82",x"20",x"25",x"D1",x"D0"
		,x"03",x"4C",x"20",x"E1",x"A5",x"83",x"C9",x"0F"
		,x"F0",x"5A",x"B5",x"F2",x"29",x"08",x"D0",x"13"
		,x"20",x"25",x"D1",x"C9",x"07",x"D0",x"07",x"A9"
		,x"89",x"95",x"F2",x"4C",x"DE",x"D3",x"A9",x"00"
		,x"95",x"F2",x"60",x"A5",x"83",x"F0",x"32",x"20"
		,x"25",x"D1",x"C9",x"04",x"90",x"22",x"20",x"2F"
		,x"D1",x"B5",x"99",x"D9",x"44",x"02",x"D0",x"04"
		,x"A9",x"00",x"95",x"99",x"F6",x"99",x"A1",x"99"
		,x"99",x"3E",x"02",x"B5",x"99",x"D9",x"44",x"02"
		,x"D0",x"05",x"A9",x"81",x"99",x"F2",x"00",x"60"
		,x"20",x"56",x"D1",x"A6",x"82",x"9D",x"3E",x"02"
		,x"60",x"AD",x"54",x"02",x"F0",x"F2",x"20",x"67"
		,x"ED",x"4C",x"03",x"D4",x"20",x"E8",x"D4",x"C9"
		,x"D4",x"D0",x"18",x"A5",x"95",x"C9",x"02",x"D0"
		,x"12",x"A9",x"0D",x"85",x"85",x"20",x"23",x"C1"
		,x"A9",x"00",x"20",x"C1",x"E6",x"C6",x"A5",x"A9"
		,x"80",x"D0",x"12",x"20",x"37",x"D1",x"85",x"85"
		,x"D0",x"09",x"A9",x"D4",x"20",x"C8",x"D4",x"A9"
		,x"02",x"95",x"9A",x"A9",x"88",x"85",x"F7",x"A5"
		,x"85",x"8D",x"43",x"02",x"60",x"20",x"93",x"DF"
		,x"0A",x"AA",x"A9",x"00",x"95",x"99",x"A1",x"99"
		,x"F0",x"05",x"D6",x"99",x"4C",x"56",x"D1",x"60"
		,x"A9",x"80",x"D0",x"02",x"A9",x"90",x"05",x"7F"
		,x"8D",x"4D",x"02",x"A5",x"F9",x"20",x"D3",x"D6"
		,x"A6",x"F9",x"4C",x"93",x"D5",x"A9",x"01",x"8D"
		,x"4A",x"02",x"A9",x"11",x"85",x"83",x"20",x"46"
		,x"DC",x"A9",x"02",x"4C",x"C8",x"D4",x"A9",x"12"
		,x"85",x"83",x"4C",x"DA",x"DC",x"20",x"3B",x"DE"
		,x"A9",x"01",x"85",x"6F",x"A5",x"69",x"48",x"A9"
		,x"03",x"85",x"69",x"20",x"2D",x"F1",x"68",x"85"
		,x"69",x"A9",x"00",x"20",x"C8",x"D4",x"A5",x"80"
		,x"20",x"F1",x"CF",x"A5",x"81",x"20",x"F1",x"CF"
		,x"20",x"C7",x"D0",x"20",x"99",x"D5",x"A9",x"00"
		,x"20",x"C8",x"D4",x"20",x"F1",x"CF",x"D0",x"FB"
		,x"20",x"F1",x"CF",x"A9",x"FF",x"4C",x"F1",x"CF"
		,x"85",x"6F",x"20",x"93",x"DF",x"0A",x"AA",x"B5"
		,x"9A",x"85",x"95",x"A5",x"6F",x"95",x"99",x"85"
		,x"94",x"60",x"A9",x"11",x"85",x"83",x"20",x"27"
		,x"D2",x"A9",x"12",x"85",x"83",x"4C",x"27",x"D2"
		,x"20",x"93",x"DF",x"0A",x"AA",x"B5",x"9A",x"85"
		,x"95",x"B5",x"99",x"85",x"94",x"60",x"85",x"71"
		,x"20",x"93",x"DF",x"AA",x"BD",x"E0",x"FE",x"85"
		,x"72",x"A0",x"00",x"B1",x"71",x"60",x"BD",x"5B"
		,x"02",x"29",x"01",x"0D",x"4D",x"02",x"48",x"86"
		,x"F9",x"8A",x"0A",x"AA",x"B5",x"07",x"8D",x"4D"
		,x"02",x"B5",x"06",x"F0",x"2D",x"CD",x"D7",x"FE"
		,x"B0",x"28",x"AA",x"68",x"48",x"29",x"F0",x"C9"
		,x"90",x"D0",x"4F",x"68",x"48",x"4A",x"B0",x"05"
		,x"AD",x"01",x"01",x"90",x"03",x"AD",x"02",x"01"
		,x"F0",x"05",x"CD",x"D5",x"FE",x"D0",x"33",x"8A"
		,x"20",x"4B",x"F2",x"CD",x"4D",x"02",x"F0",x"02"
		,x"B0",x"30",x"20",x"52",x"D5",x"A9",x"66",x"4C"
		,x"45",x"E6",x"A5",x"F9",x"0A",x"AA",x"B5",x"06"
		,x"85",x"80",x"B5",x"07",x"85",x"81",x"60",x"A5"
		,x"80",x"F0",x"EA",x"CD",x"D7",x"FE",x"B0",x"E5"
		,x"20",x"4B",x"F2",x"C5",x"81",x"F0",x"DE",x"90"
		,x"DC",x"60",x"20",x"52",x"D5",x"A9",x"73",x"4C"
		,x"45",x"E6",x"A6",x"F9",x"68",x"8D",x"4D",x"02"
		,x"95",x"00",x"9D",x"5B",x"02",x"60",x"A9",x"80"
		,x"D0",x"02",x"A9",x"90",x"05",x"7F",x"A6",x"F9"
		,x"8D",x"4D",x"02",x"AD",x"4D",x"02",x"20",x"0E"
		,x"D5",x"20",x"A6",x"D5",x"B0",x"FB",x"48",x"A9"
		,x"00",x"8D",x"98",x"02",x"68",x"60",x"B5",x"00"
		,x"30",x"1A",x"C9",x"02",x"90",x"14",x"C9",x"08"
		,x"F0",x"08",x"C9",x"0B",x"F0",x"04",x"C9",x"0F"
		,x"D0",x"0C",x"2C",x"98",x"02",x"30",x"03",x"4C"
		,x"3F",x"D6",x"18",x"60",x"38",x"60",x"98",x"48"
		,x"A5",x"7F",x"48",x"BD",x"5B",x"02",x"29",x"01"
		,x"85",x"7F",x"A8",x"B9",x"CA",x"FE",x"8D",x"6D"
		,x"02",x"20",x"A6",x"D6",x"C9",x"02",x"B0",x"03"
		,x"4C",x"6D",x"D6",x"BD",x"5B",x"02",x"29",x"F0"
		,x"48",x"C9",x"90",x"D0",x"07",x"A5",x"7F",x"09"
		,x"B8",x"9D",x"5B",x"02",x"24",x"6A",x"70",x"39"
		,x"A9",x"00",x"8D",x"99",x"02",x"8D",x"9A",x"02"
		,x"AC",x"99",x"02",x"AD",x"9A",x"02",x"38",x"F9"
		,x"DB",x"FE",x"8D",x"9A",x"02",x"B9",x"DB",x"FE"
		,x"20",x"76",x"D6",x"EE",x"99",x"02",x"20",x"A6"
		,x"D6",x"C9",x"02",x"90",x"08",x"AC",x"99",x"02"
		,x"B9",x"DB",x"FE",x"D0",x"DB",x"AD",x"9A",x"02"
		,x"20",x"76",x"D6",x"B5",x"00",x"C9",x"02",x"90"
		,x"2B",x"24",x"6A",x"10",x"0F",x"68",x"C9",x"90"
		,x"D0",x"05",x"05",x"7F",x"9D",x"5B",x"02",x"B5"
		,x"00",x"20",x"0A",x"E6",x"68",x"2C",x"98",x"02"
		,x"30",x"23",x"48",x"A9",x"C0",x"05",x"7F",x"95"
		,x"00",x"B5",x"00",x"30",x"FC",x"20",x"A6",x"D6"
		,x"C9",x"02",x"B0",x"D9",x"68",x"C9",x"90",x"D0"
		,x"0C",x"05",x"7F",x"9D",x"5B",x"02",x"20",x"A6"
		,x"D6",x"C9",x"02",x"B0",x"D2",x"68",x"85",x"7F"
		,x"68",x"A8",x"B5",x"00",x"18",x"60",x"C9",x"00"
		,x"F0",x"18",x"30",x"0C",x"A0",x"01",x"20",x"93"
		,x"D6",x"38",x"E9",x"01",x"D0",x"F6",x"F0",x"0A"
		,x"A0",x"FF",x"20",x"93",x"D6",x"18",x"69",x"01"
		,x"D0",x"F6",x"60",x"48",x"98",x"A4",x"7F",x"99"
		,x"FE",x"02",x"D9",x"FE",x"02",x"F0",x"FB",x"A9"
		,x"00",x"99",x"FE",x"02",x"68",x"60",x"A5",x"6A"
		,x"29",x"3F",x"A8",x"AD",x"6D",x"02",x"4D",x"00"
		,x"1C",x"8D",x"00",x"1C",x"BD",x"5B",x"02",x"95"
		,x"00",x"B5",x"00",x"30",x"FC",x"C9",x"02",x"90"
		,x"03",x"88",x"D0",x"E7",x"48",x"AD",x"6D",x"02"
		,x"0D",x"00",x"1C",x"8D",x"00",x"1C",x"68",x"60"
		,x"20",x"93",x"DF",x"0A",x"A8",x"A5",x"80",x"99"
		,x"06",x"00",x"A5",x"81",x"99",x"07",x"00",x"A5"
		,x"7F",x"0A",x"AA",x"60",x"A5",x"83",x"48",x"A5"
		,x"82",x"48",x"A5",x"81",x"48",x"A5",x"80",x"48"
		,x"A9",x"11",x"85",x"83",x"20",x"3B",x"DE",x"AD"
		,x"4A",x"02",x"48",x"A5",x"E2",x"29",x"01",x"85"
		,x"7F",x"A6",x"F9",x"5D",x"5B",x"02",x"4A",x"90"
		,x"0C",x"A2",x"01",x"8E",x"92",x"02",x"20",x"AC"
		,x"C5",x"F0",x"1D",x"D0",x"28",x"AD",x"91",x"02"
		,x"F0",x"0C",x"C5",x"81",x"F0",x"1F",x"85",x"81"
		,x"20",x"60",x"D4",x"4C",x"3D",x"D7",x"A9",x"01"
		,x"8D",x"92",x"02",x"20",x"17",x"C6",x"D0",x"0D"
		,x"20",x"8D",x"D4",x"A5",x"81",x"8D",x"91",x"02"
		,x"A9",x"02",x"8D",x"92",x"02",x"AD",x"92",x"02"
		,x"20",x"C8",x"D4",x"68",x"8D",x"4A",x"02",x"C9"
		,x"04",x"D0",x"02",x"09",x"80",x"20",x"F1",x"CF"
		,x"68",x"8D",x"80",x"02",x"20",x"F1",x"CF",x"68"
		,x"8D",x"85",x"02",x"20",x"F1",x"CF",x"20",x"93"
		,x"DF",x"A8",x"AD",x"7A",x"02",x"AA",x"A9",x"10"
		,x"20",x"6E",x"C6",x"A0",x"10",x"A9",x"00",x"91"
		,x"94",x"C8",x"C0",x"1B",x"90",x"F9",x"AD",x"4A"
		,x"02",x"C9",x"04",x"D0",x"13",x"A0",x"10",x"AD"
		,x"59",x"02",x"91",x"94",x"C8",x"AD",x"5A",x"02"
		,x"91",x"94",x"C8",x"AD",x"58",x"02",x"91",x"94"
		,x"20",x"64",x"D4",x"68",x"85",x"82",x"AA",x"68"
		,x"85",x"83",x"AD",x"91",x"02",x"85",x"D8",x"9D"
		,x"60",x"02",x"AD",x"92",x"02",x"85",x"DD",x"9D"
		,x"66",x"02",x"AD",x"4A",x"02",x"85",x"E7",x"A5"
		,x"7F",x"85",x"E2",x"60",x"A5",x"83",x"8D",x"4C"
		,x"02",x"20",x"B3",x"C2",x"8E",x"2A",x"02",x"AE"
		,x"00",x"02",x"AD",x"4C",x"02",x"D0",x"2C",x"E0"
		,x"2A",x"D0",x"28",x"A5",x"7E",x"F0",x"4D",x"85"
		,x"80",x"AD",x"6E",x"02",x"85",x"7F",x"85",x"E2"
		,x"A9",x"02",x"85",x"E7",x"AD",x"6F",x"02",x"85"
		,x"81",x"20",x"00",x"C1",x"20",x"46",x"DC",x"A9"
		,x"04",x"05",x"7F",x"A6",x"82",x"99",x"EC",x"00"
		,x"4C",x"94",x"C1",x"E0",x"24",x"D0",x"1E",x"AD"
		,x"4C",x"02",x"D0",x"03",x"4C",x"55",x"DA",x"20"
		,x"D1",x"C1",x"AD",x"85",x"FE",x"85",x"80",x"A9"
		,x"00",x"85",x"81",x"20",x"46",x"DC",x"A5",x"7F"
		,x"09",x"02",x"4C",x"EB",x"D7",x"E0",x"23",x"D0"
		,x"12",x"4C",x"84",x"CB",x"A9",x"02",x"8D",x"96"
		,x"02",x"A9",x"00",x"85",x"7F",x"8D",x"8E",x"02"
		,x"20",x"42",x"D0",x"20",x"E5",x"C1",x"D0",x"04"
		,x"A2",x"00",x"F0",x"0C",x"8A",x"F0",x"05",x"A9"
		,x"30",x"4C",x"C8",x"C1",x"88",x"F0",x"01",x"88"
		,x"8C",x"7A",x"02",x"A9",x"8D",x"20",x"68",x"C2"
		,x"E8",x"8E",x"78",x"02",x"20",x"12",x"C3",x"20"
		,x"CA",x"C3",x"20",x"9D",x"C4",x"A2",x"00",x"8E"
		,x"58",x"02",x"8E",x"97",x"02",x"8E",x"4A",x"02"
		,x"E8",x"EC",x"77",x"02",x"B0",x"10",x"20",x"09"
		,x"DA",x"E8",x"EC",x"77",x"02",x"B0",x"07",x"C0"
		,x"04",x"F0",x"3E",x"20",x"09",x"DA",x"AE",x"4C"
		,x"02",x"86",x"83",x"E0",x"02",x"B0",x"12",x"8E"
		,x"97",x"02",x"A9",x"40",x"8D",x"F9",x"02",x"AD"
		,x"4A",x"02",x"D0",x"1B",x"A9",x"02",x"8D",x"4A"
		,x"02",x"AD",x"4A",x"02",x"D0",x"11",x"A5",x"E7"
		,x"29",x"07",x"8D",x"4A",x"02",x"AD",x"80",x"02"
		,x"D0",x"05",x"A9",x"01",x"8D",x"4A",x"02",x"AD"
		,x"97",x"02",x"C9",x"01",x"F0",x"18",x"4C",x"40"
		,x"D9",x"BC",x"7A",x"02",x"B9",x"00",x"02",x"8D"
		,x"58",x"02",x"AD",x"80",x"02",x"D0",x"B7",x"A9"
		,x"01",x"8D",x"97",x"02",x"D0",x"B0",x"A5",x"E7"
		,x"29",x"80",x"AA",x"D0",x"14",x"A9",x"20",x"24"
		,x"E7",x"F0",x"06",x"20",x"B6",x"C8",x"4C",x"E3"
		,x"D9",x"AD",x"80",x"02",x"D0",x"03",x"4C",x"E3"
		,x"D9",x"AD",x"00",x"02",x"C9",x"40",x"F0",x"0D"
		,x"8A",x"D0",x"05",x"A9",x"63",x"4C",x"C8",x"C1"
		,x"A9",x"33",x"4C",x"C8",x"C1",x"A5",x"E7",x"29"
		,x"07",x"CD",x"4A",x"02",x"D0",x"67",x"C9",x"04"
		,x"F0",x"63",x"20",x"DA",x"DC",x"A5",x"82",x"8D"
		,x"70",x"02",x"A9",x"11",x"85",x"83",x"20",x"EB"
		,x"D0",x"AD",x"94",x"02",x"20",x"C8",x"D4",x"A0"
		,x"00",x"B1",x"94",x"09",x"20",x"91",x"94",x"A0"
		,x"1A",x"A5",x"80",x"91",x"94",x"C8",x"A5",x"81"
		,x"91",x"94",x"AE",x"70",x"02",x"A5",x"D8",x"9D"
		,x"60",x"02",x"A5",x"DD",x"9D",x"66",x"02",x"20"
		,x"3B",x"DE",x"20",x"64",x"D4",x"4C",x"EF",x"D9"
		,x"AD",x"80",x"02",x"D0",x"05",x"A9",x"62",x"4C"
		,x"C8",x"C1",x"AD",x"97",x"02",x"C9",x"03",x"F0"
		,x"0B",x"A9",x"20",x"24",x"E7",x"F0",x"05",x"A9"
		,x"60",x"4C",x"C8",x"C1",x"A5",x"E7",x"29",x"07"
		,x"CD",x"4A",x"02",x"F0",x"05",x"A9",x"64",x"4C"
		,x"C8",x"C1",x"A0",x"00",x"8C",x"79",x"02",x"AE"
		,x"97",x"02",x"E0",x"02",x"D0",x"1A",x"C9",x"04"
		,x"F0",x"EB",x"B1",x"94",x"29",x"4F",x"91",x"94"
		,x"A5",x"83",x"48",x"A9",x"11",x"85",x"83",x"20"
		,x"3B",x"DE",x"20",x"64",x"D4",x"68",x"85",x"83"
		,x"20",x"A0",x"D9",x"AD",x"97",x"02",x"C9",x"02"
		,x"D0",x"55",x"20",x"2A",x"DA",x"4C",x"94",x"C1"
		,x"A0",x"13",x"B1",x"94",x"8D",x"59",x"02",x"C8"
		,x"B1",x"94",x"8D",x"5A",x"02",x"C8",x"B1",x"94"
		,x"AE",x"58",x"02",x"8D",x"58",x"02",x"8A",x"F0"
		,x"0A",x"CD",x"58",x"02",x"F0",x"05",x"A9",x"50"
		,x"20",x"C8",x"C1",x"AE",x"79",x"02",x"BD",x"80"
		,x"02",x"85",x"80",x"BD",x"85",x"02",x"85",x"81"
		,x"20",x"46",x"DC",x"A4",x"82",x"AE",x"79",x"02"
		,x"B5",x"D8",x"99",x"60",x"02",x"B5",x"DD",x"99"
		,x"66",x"02",x"60",x"A5",x"E2",x"29",x"01",x"85"
		,x"7F",x"20",x"DA",x"DC",x"20",x"E4",x"D6",x"A5"
		,x"83",x"C9",x"02",x"B0",x"11",x"20",x"3E",x"DE"
		,x"A5",x"80",x"85",x"7E",x"A5",x"7F",x"8D",x"6E"
		,x"02",x"A5",x"81",x"8D",x"6F",x"02",x"4C",x"99"
		,x"C1",x"BC",x"7A",x"02",x"B9",x"00",x"02",x"A0"
		,x"04",x"88",x"30",x"08",x"D9",x"B2",x"FE",x"D0"
		,x"F8",x"8C",x"97",x"02",x"A0",x"05",x"88",x"30"
		,x"08",x"D9",x"B6",x"FE",x"D0",x"F8",x"8C",x"4A"
		,x"02",x"60",x"20",x"39",x"CA",x"A9",x"80",x"20"
		,x"A6",x"DD",x"F0",x"F6",x"20",x"95",x"DE",x"A6"
		,x"81",x"E8",x"8A",x"D0",x"05",x"20",x"A3",x"D1"
		,x"A9",x"02",x"20",x"C8",x"D4",x"A6",x"82",x"A9"
		,x"01",x"95",x"F2",x"A9",x"80",x"05",x"82",x"A6"
		,x"83",x"9D",x"2B",x"02",x"60",x"A9",x"0C",x"8D"
		,x"2A",x"02",x"A9",x"00",x"AE",x"74",x"02",x"CA"
		,x"F0",x"0B",x"CA",x"D0",x"21",x"AD",x"01",x"02"
		,x"20",x"BD",x"C3",x"30",x"19",x"85",x"E2",x"EE"
		,x"77",x"02",x"EE",x"78",x"02",x"EE",x"7A",x"02"
		,x"A9",x"80",x"85",x"E7",x"A9",x"2A",x"8D",x"00"
		,x"02",x"8D",x"01",x"02",x"D0",x"18",x"20",x"E5"
		,x"C1",x"D0",x"05",x"20",x"DC",x"C2",x"A0",x"03"
		,x"88",x"88",x"8C",x"7A",x"02",x"20",x"00",x"C2"
		,x"20",x"98",x"C3",x"20",x"20",x"C3",x"20",x"CA"
		,x"C3",x"20",x"B7",x"C7",x"20",x"9D",x"C4",x"20"
		,x"9E",x"EC",x"20",x"37",x"D1",x"A6",x"82",x"9D"
		,x"3E",x"02",x"A5",x"7F",x"8D",x"8E",x"02",x"09"
		,x"04",x"95",x"EC",x"A9",x"00",x"85",x"A3",x"60"
		,x"A9",x"00",x"8D",x"F9",x"02",x"A5",x"83",x"D0"
		,x"0B",x"A9",x"00",x"8D",x"54",x"02",x"20",x"27"
		,x"D2",x"4C",x"DA",x"D4",x"C9",x"0F",x"F0",x"14"
		,x"20",x"02",x"DB",x"A5",x"83",x"C9",x"02",x"90"
		,x"F0",x"AD",x"6C",x"02",x"D0",x"03",x"4C",x"94"
		,x"C1",x"4C",x"AD",x"C1",x"A9",x"0E",x"85",x"83"
		,x"20",x"02",x"DB",x"C6",x"83",x"10",x"F9",x"AD"
		,x"6C",x"02",x"D0",x"03",x"4C",x"94",x"C1",x"4C"
		,x"AD",x"C1",x"A6",x"83",x"BD",x"2B",x"02",x"C9"
		,x"FF",x"D0",x"01",x"60",x"29",x"0F",x"85",x"82"
		,x"20",x"25",x"D1",x"C9",x"07",x"F0",x"0F",x"C9"
		,x"04",x"F0",x"11",x"20",x"07",x"D1",x"B0",x"09"
		,x"20",x"62",x"DB",x"20",x"A5",x"DB",x"20",x"F4"
		,x"EE",x"4C",x"27",x"D2",x"20",x"F1",x"DD",x"20"
		,x"1E",x"CF",x"20",x"CB",x"E1",x"A6",x"D5",x"86"
		,x"73",x"E6",x"73",x"A9",x"00",x"85",x"70",x"85"
		,x"71",x"A5",x"D6",x"38",x"E9",x"0E",x"85",x"72"
		,x"20",x"51",x"DF",x"A6",x"82",x"A5",x"70",x"95"
		,x"B5",x"A5",x"71",x"95",x"BB",x"A9",x"40",x"20"
		,x"A6",x"DD",x"F0",x"03",x"20",x"A5",x"DB",x"4C"
		,x"27",x"D2",x"A6",x"82",x"B5",x"B5",x"15",x"BB"
		,x"D0",x"0C",x"20",x"E8",x"D4",x"C9",x"02",x"D0"
		,x"05",x"A9",x"0D",x"20",x"F1",x"CF",x"20",x"E8"
		,x"D4",x"C9",x"02",x"D0",x"0F",x"20",x"1E",x"CF"
		,x"A6",x"82",x"B5",x"B5",x"D0",x"02",x"D6",x"BB"
		,x"D6",x"B5",x"A9",x"00",x"38",x"E9",x"01",x"48"
		,x"A9",x"00",x"20",x"C8",x"D4",x"20",x"F1",x"CF"
		,x"68",x"20",x"F1",x"CF",x"20",x"C7",x"D0",x"20"
		,x"99",x"D5",x"4C",x"1E",x"CF",x"A6",x"82",x"8E"
		,x"70",x"02",x"A5",x"83",x"48",x"BD",x"60",x"02"
		,x"85",x"81",x"BD",x"66",x"02",x"8D",x"94",x"02"
		,x"B5",x"EC",x"29",x"01",x"85",x"7F",x"AD",x"85"
		,x"FE",x"85",x"80",x"20",x"93",x"DF",x"48",x"85"
		,x"F9",x"20",x"60",x"D4",x"A0",x"00",x"BD",x"E0"
		,x"FE",x"85",x"87",x"AD",x"94",x"02",x"85",x"86"
		,x"B1",x"86",x"29",x"20",x"F0",x"43",x"20",x"25"
		,x"D1",x"C9",x"04",x"F0",x"44",x"B1",x"86",x"29"
		,x"8F",x"91",x"86",x"C8",x"B1",x"86",x"85",x"80"
		,x"84",x"71",x"A0",x"1B",x"B1",x"86",x"48",x"88"
		,x"B1",x"86",x"D0",x"0A",x"85",x"80",x"68",x"85"
		,x"81",x"A9",x"67",x"20",x"45",x"E6",x"48",x"A9"
		,x"00",x"91",x"86",x"C8",x"91",x"86",x"68",x"A4"
		,x"71",x"91",x"86",x"C8",x"B1",x"86",x"85",x"81"
		,x"68",x"91",x"86",x"20",x"7D",x"C8",x"4C",x"29"
		,x"DC",x"B1",x"86",x"29",x"0F",x"09",x"80",x"91"
		,x"86",x"AE",x"70",x"02",x"A0",x"1C",x"B5",x"B5"
		,x"91",x"86",x"C8",x"B5",x"BB",x"91",x"86",x"68"
		,x"AA",x"A9",x"90",x"05",x"7F",x"20",x"90",x"D5"
		,x"68",x"85",x"83",x"4C",x"07",x"D1",x"A9",x"01"
		,x"20",x"E2",x"D1",x"20",x"B6",x"DC",x"AD",x"4A"
		,x"02",x"48",x"0A",x"05",x"7F",x"95",x"EC",x"20"
		,x"9B",x"D0",x"A6",x"82",x"A5",x"80",x"D0",x"05"
		,x"A5",x"81",x"9D",x"44",x"02",x"68",x"C9",x"04"
		,x"D0",x"3F",x"A4",x"83",x"B9",x"2B",x"02",x"09"
		,x"40",x"99",x"2B",x"02",x"AD",x"58",x"02",x"95"
		,x"C7",x"20",x"8E",x"D2",x"10",x"03",x"4C",x"0F"
		,x"D2",x"A6",x"82",x"95",x"CD",x"AC",x"59",x"02"
		,x"84",x"80",x"AC",x"5A",x"02",x"84",x"81",x"20"
		,x"D3",x"D6",x"20",x"73",x"DE",x"20",x"99",x"D5"
		,x"A6",x"82",x"A9",x"02",x"95",x"C1",x"A9",x"00"
		,x"20",x"C8",x"D4",x"20",x"53",x"E1",x"4C",x"3E"
		,x"DE",x"20",x"56",x"D1",x"A6",x"82",x"9D",x"3E"
		,x"02",x"A9",x"88",x"95",x"F2",x"60",x"A6",x"82"
		,x"B5",x"A7",x"0A",x"30",x"06",x"A8",x"A9",x"02"
		,x"99",x"99",x"00",x"B5",x"AE",x"09",x"80",x"95"
		,x"AE",x"0A",x"30",x"06",x"A8",x"A9",x"02",x"99"
		,x"99",x"00",x"A9",x"00",x"95",x"B5",x"4C",x"75"
		,x"C0",x"EA",x"20",x"A9",x"F1",x"A9",x"01",x"20"
		,x"DF",x"D1",x"20",x"D0",x"D6",x"20",x"B6",x"DC"
		,x"A6",x"82",x"AD",x"4A",x"02",x"48",x"0A",x"05"
		,x"7F",x"95",x"EC",x"68",x"C9",x"04",x"F0",x"05"
		,x"A9",x"01",x"95",x"F2",x"60",x"A4",x"83",x"B9"
		,x"2B",x"02",x"29",x"3F",x"09",x"40",x"99",x"2B"
		,x"02",x"AD",x"58",x"02",x"95",x"C7",x"20",x"8E"
		,x"D2",x"10",x"03",x"4C",x"0F",x"D2",x"A6",x"82"
		,x"95",x"CD",x"20",x"C1",x"DE",x"20",x"1E",x"F1"
		,x"A5",x"80",x"8D",x"59",x"02",x"A5",x"81",x"8D"
		,x"5A",x"02",x"A6",x"82",x"B5",x"CD",x"20",x"D3"
		,x"D6",x"A9",x"00",x"20",x"E9",x"DE",x"A9",x"00"
		,x"20",x"8D",x"DD",x"A9",x"11",x"20",x"8D",x"DD"
		,x"A9",x"00",x"20",x"8D",x"DD",x"AD",x"58",x"02"
		,x"20",x"8D",x"DD",x"A5",x"80",x"20",x"8D",x"DD"
		,x"A5",x"81",x"20",x"8D",x"DD",x"A9",x"10",x"20"
		,x"E9",x"DE",x"20",x"3E",x"DE",x"A5",x"80",x"20"
		,x"8D",x"DD",x"A5",x"81",x"20",x"8D",x"DD",x"20"
		,x"6C",x"DE",x"20",x"99",x"D5",x"A9",x"02",x"20"
		,x"C8",x"D4",x"A6",x"82",x"38",x"A9",x"00",x"F5"
		,x"C7",x"95",x"C1",x"20",x"E2",x"E2",x"20",x"19"
		,x"DE",x"20",x"5E",x"DE",x"20",x"99",x"D5",x"20"
		,x"F4",x"EE",x"4C",x"98",x"DC",x"48",x"A6",x"82"
		,x"B5",x"CD",x"4C",x"FD",x"CF",x"90",x"06",x"A6"
		,x"82",x"15",x"EC",x"D0",x"06",x"A6",x"82",x"49"
		,x"FF",x"35",x"EC",x"95",x"EC",x"60",x"A6",x"82"
		,x"35",x"EC",x"60",x"20",x"93",x"DF",x"AA",x"BD"
		,x"5B",x"02",x"29",x"F0",x"C9",x"90",x"60",x"A2"
		,x"00",x"86",x"71",x"BD",x"2B",x"02",x"C9",x"FF"
		,x"D0",x"08",x"A6",x"71",x"E8",x"E0",x"10",x"90"
		,x"F0",x"60",x"86",x"71",x"29",x"3F",x"A8",x"B9"
		,x"EC",x"00",x"29",x"01",x"85",x"70",x"AE",x"53"
		,x"02",x"B5",x"E2",x"29",x"01",x"C5",x"70",x"D0"
		,x"E1",x"B9",x"60",x"02",x"D5",x"D8",x"D0",x"DA"
		,x"B9",x"66",x"02",x"D5",x"DD",x"D0",x"D3",x"18"
		,x"60",x"20",x"9E",x"DF",x"50",x"06",x"20",x"5E"
		,x"DE",x"20",x"99",x"D5",x"60",x"20",x"2B",x"DE"
		,x"A5",x"80",x"91",x"94",x"C8",x"A5",x"81",x"91"
		,x"94",x"4C",x"05",x"E1",x"20",x"2B",x"DE",x"B1"
		,x"94",x"85",x"80",x"C8",x"B1",x"94",x"85",x"81"
		,x"60",x"20",x"2B",x"DE",x"A9",x"00",x"91",x"94"
		,x"C8",x"A6",x"82",x"B5",x"C1",x"AA",x"CA",x"8A"
		,x"91",x"94",x"60",x"20",x"93",x"DF",x"0A",x"AA"
		,x"B5",x"9A",x"85",x"95",x"A9",x"00",x"85",x"94"
		,x"A0",x"00",x"60",x"20",x"EB",x"D0",x"20",x"93"
		,x"DF",x"85",x"F9",x"0A",x"A8",x"B9",x"06",x"00"
		,x"85",x"80",x"B9",x"07",x"00",x"85",x"81",x"60"
		,x"A9",x"90",x"8D",x"4D",x"02",x"D0",x"28",x"A9"
		,x"80",x"8D",x"4D",x"02",x"D0",x"21",x"A9",x"90"
		,x"8D",x"4D",x"02",x"D0",x"26",x"A9",x"80",x"8D"
		,x"4D",x"02",x"D0",x"1F",x"A9",x"90",x"8D",x"4D"
		,x"02",x"D0",x"02",x"A9",x"80",x"8D",x"4D",x"02"
		,x"A6",x"82",x"B5",x"CD",x"AA",x"10",x"13",x"20"
		,x"D0",x"D6",x"20",x"93",x"DF",x"AA",x"A5",x"7F"
		,x"9D",x"5B",x"02",x"20",x"15",x"E1",x"20",x"93"
		,x"DF",x"AA",x"4C",x"06",x"D5",x"A9",x"00",x"20"
		,x"C8",x"D4",x"20",x"37",x"D1",x"85",x"80",x"20"
		,x"37",x"D1",x"85",x"81",x"60",x"48",x"A9",x"00"
		,x"85",x"6F",x"85",x"71",x"B9",x"E0",x"FE",x"85"
		,x"70",x"BD",x"E0",x"FE",x"85",x"72",x"68",x"A8"
		,x"88",x"B1",x"6F",x"91",x"71",x"88",x"10",x"F9"
		,x"60",x"A8",x"B9",x"E0",x"FE",x"85",x"70",x"A9"
		,x"00",x"85",x"6F",x"A8",x"91",x"6F",x"C8",x"D0"
		,x"FB",x"60",x"A9",x"00",x"20",x"DC",x"DE",x"A0"
		,x"02",x"B1",x"94",x"60",x"85",x"94",x"A6",x"82"
		,x"B5",x"CD",x"AA",x"BD",x"E0",x"FE",x"85",x"95"
		,x"60",x"48",x"20",x"DC",x"DE",x"48",x"8A",x"0A"
		,x"AA",x"68",x"95",x"9A",x"68",x"95",x"99",x"60"
		,x"20",x"66",x"DF",x"30",x"0E",x"50",x"13",x"A6"
		,x"82",x"B5",x"CD",x"20",x"1B",x"DF",x"20",x"66"
		,x"DF",x"10",x"07",x"20",x"CB",x"E1",x"2C",x"CE"
		,x"FE",x"60",x"A5",x"D6",x"20",x"E9",x"DE",x"2C"
		,x"CD",x"FE",x"60",x"85",x"F9",x"A9",x"80",x"D0"
		,x"04",x"85",x"F9",x"A9",x"90",x"48",x"B5",x"EC"
		,x"29",x"01",x"85",x"7F",x"68",x"05",x"7F",x"8D"
		,x"4D",x"02",x"B1",x"94",x"85",x"80",x"C8",x"B1"
		,x"94",x"85",x"81",x"A5",x"F9",x"20",x"D3",x"D6"
		,x"A6",x"F9",x"4C",x"93",x"D5",x"A6",x"82",x"B5"
		,x"CD",x"4C",x"EB",x"D4",x"A9",x"78",x"20",x"5C"
		,x"DF",x"CA",x"10",x"F8",x"A5",x"72",x"4A",x"20"
		,x"5C",x"DF",x"A5",x"73",x"18",x"65",x"70",x"85"
		,x"70",x"90",x"02",x"E6",x"71",x"60",x"20",x"D2"
		,x"DE",x"C5",x"D5",x"D0",x"0E",x"A4",x"D6",x"B1"
		,x"94",x"F0",x"04",x"2C",x"CD",x"FE",x"60",x"2C"
		,x"CF",x"FE",x"60",x"A5",x"D5",x"C9",x"06",x"B0"
		,x"0A",x"0A",x"A8",x"A9",x"04",x"85",x"94",x"B1"
		,x"94",x"D0",x"04",x"2C",x"D0",x"FE",x"60",x"2C"
		,x"CE",x"FE",x"60",x"A6",x"82",x"B5",x"A7",x"10"
		,x"02",x"B5",x"AE",x"29",x"BF",x"60",x"A6",x"82"
		,x"8E",x"57",x"02",x"B5",x"A7",x"10",x"09",x"8A"
		,x"18",x"69",x"07",x"8D",x"57",x"02",x"B5",x"AE"
		,x"85",x"70",x"29",x"1F",x"24",x"70",x"60",x"A6"
		,x"82",x"B5",x"A7",x"30",x"02",x"B5",x"AE",x"C9"
		,x"FF",x"60",x"A6",x"82",x"09",x"80",x"B4",x"A7"
		,x"10",x"03",x"95",x"A7",x"60",x"95",x"AE",x"60"
		,x"A9",x"20",x"20",x"9D",x"DD",x"A9",x"80",x"20"
		,x"A6",x"DD",x"D0",x"41",x"A6",x"82",x"F6",x"B5"
		,x"D0",x"02",x"F6",x"BB",x"A6",x"82",x"B5",x"C1"
		,x"F0",x"2E",x"20",x"E8",x"D4",x"A6",x"82",x"D5"
		,x"C1",x"90",x"03",x"20",x"3C",x"E0",x"A6",x"82"
		,x"B5",x"C1",x"20",x"C8",x"D4",x"A1",x"99",x"85"
		,x"85",x"A9",x"20",x"20",x"9D",x"DD",x"20",x"04"
		,x"E3",x"48",x"90",x"28",x"A9",x"00",x"20",x"F6"
		,x"D4",x"D0",x"21",x"68",x"C9",x"02",x"F0",x"12"
		,x"A9",x"80",x"20",x"97",x"DD",x"20",x"2F",x"D1"
		,x"B5",x"99",x"99",x"44",x"02",x"A9",x"0D",x"85"
		,x"85",x"60",x"20",x"35",x"E0",x"A6",x"82",x"A9"
		,x"00",x"95",x"C1",x"60",x"68",x"A6",x"82",x"95"
		,x"C1",x"4C",x"6E",x"E1",x"20",x"D3",x"D1",x"20"
		,x"95",x"DE",x"20",x"9E",x"DF",x"50",x"16",x"20"
		,x"5E",x"DE",x"20",x"1E",x"CF",x"A9",x"02",x"20"
		,x"C8",x"D4",x"20",x"AB",x"DD",x"D0",x"24",x"20"
		,x"57",x"DE",x"4C",x"99",x"D5",x"20",x"1E",x"CF"
		,x"20",x"AB",x"DD",x"D0",x"06",x"20",x"57",x"DE"
		,x"20",x"99",x"D5",x"20",x"95",x"DE",x"A5",x"80"
		,x"F0",x"09",x"20",x"1E",x"CF",x"20",x"57",x"DE"
		,x"20",x"1E",x"CF",x"60",x"20",x"05",x"E1",x"20"
		,x"93",x"DF",x"0A",x"AA",x"A5",x"85",x"81",x"99"
		,x"B4",x"99",x"C8",x"D0",x"09",x"A4",x"82",x"B9"
		,x"C1",x"00",x"F0",x"0A",x"A0",x"02",x"98",x"A4"
		,x"82",x"D9",x"C1",x"00",x"D0",x"05",x"A9",x"20"
		,x"4C",x"97",x"DD",x"F6",x"99",x"D0",x"03",x"20"
		,x"3C",x"E0",x"60",x"A9",x"A0",x"20",x"A6",x"DD"
		,x"D0",x"27",x"A5",x"85",x"20",x"7C",x"E0",x"A5"
		,x"F8",x"F0",x"0D",x"60",x"A9",x"20",x"20",x"A6"
		,x"DD",x"F0",x"05",x"A9",x"51",x"8D",x"6C",x"02"
		,x"20",x"F3",x"E0",x"20",x"53",x"E1",x"AD",x"6C"
		,x"02",x"F0",x"03",x"4C",x"C8",x"C1",x"4C",x"BC"
		,x"E6",x"29",x"80",x"D0",x"05",x"A5",x"F8",x"F0"
		,x"DB",x"60",x"A5",x"85",x"48",x"20",x"1C",x"E3"
		,x"68",x"85",x"85",x"A9",x"80",x"20",x"9D",x"DD"
		,x"4C",x"B2",x"E0",x"A9",x"20",x"20",x"A6",x"DD"
		,x"D0",x"0A",x"A9",x"00",x"85",x"85",x"20",x"7C"
		,x"E0",x"4C",x"F3",x"E0",x"60",x"A9",x"40",x"20"
		,x"97",x"DD",x"20",x"9E",x"DF",x"09",x"40",x"AE"
		,x"57",x"02",x"95",x"A7",x"60",x"20",x"9E",x"DF"
		,x"29",x"BF",x"AE",x"57",x"02",x"95",x"A7",x"60"
		,x"A9",x"80",x"20",x"A6",x"DD",x"D0",x"37",x"20"
		,x"2F",x"D1",x"B5",x"99",x"D9",x"44",x"02",x"F0"
		,x"22",x"F6",x"99",x"D0",x"06",x"20",x"3C",x"E0"
		,x"20",x"2F",x"D1",x"A1",x"99",x"99",x"3E",x"02"
		,x"A9",x"89",x"99",x"F2",x"00",x"B5",x"99",x"D9"
		,x"44",x"02",x"F0",x"01",x"60",x"A9",x"81",x"99"
		,x"F2",x"00",x"60",x"20",x"D0",x"DF",x"20",x"2F"
		,x"D1",x"A5",x"85",x"4C",x"3D",x"E1",x"A6",x"82"
		,x"A9",x"0D",x"9D",x"3E",x"02",x"A9",x"81",x"95"
		,x"F2",x"A9",x"50",x"20",x"C8",x"C1",x"A6",x"82"
		,x"B5",x"C1",x"85",x"87",x"C6",x"87",x"C9",x"02"
		,x"D0",x"04",x"A9",x"FF",x"85",x"87",x"B5",x"C7"
		,x"85",x"88",x"20",x"E8",x"D4",x"A6",x"82",x"C5"
		,x"87",x"90",x"19",x"F0",x"17",x"20",x"1E",x"CF"
		,x"20",x"B2",x"E1",x"90",x"08",x"A6",x"82",x"9D"
		,x"44",x"02",x"4C",x"1E",x"CF",x"20",x"1E",x"CF"
		,x"A9",x"FF",x"85",x"87",x"20",x"B2",x"E1",x"B0"
		,x"03",x"20",x"E8",x"D4",x"A6",x"82",x"9D",x"44"
		,x"02",x"60",x"20",x"2B",x"DE",x"A4",x"87",x"B1"
		,x"94",x"D0",x"0D",x"88",x"C0",x"02",x"90",x"04"
		,x"C6",x"88",x"D0",x"F3",x"C6",x"88",x"18",x"60"
		,x"98",x"38",x"60",x"20",x"D2",x"DE",x"85",x"D5"
		,x"A9",x"04",x"85",x"94",x"A0",x"0A",x"D0",x"04"
		,x"88",x"88",x"30",x"26",x"B1",x"94",x"F0",x"F8"
		,x"98",x"4A",x"C5",x"D5",x"F0",x"09",x"85",x"D5"
		,x"A6",x"82",x"B5",x"CD",x"20",x"1B",x"DF",x"A0"
		,x"00",x"84",x"94",x"B1",x"94",x"D0",x"0B",x"C8"
		,x"B1",x"94",x"A8",x"88",x"84",x"D6",x"98",x"4C"
		,x"E9",x"DE",x"A9",x"67",x"20",x"45",x"E6",x"20"
		,x"B3",x"C2",x"AD",x"01",x"02",x"85",x"83",x"20"
		,x"EB",x"D0",x"90",x"05",x"A9",x"70",x"20",x"C8"
		,x"C1",x"A9",x"A0",x"20",x"9D",x"DD",x"20",x"25"
		,x"D1",x"F0",x"05",x"A9",x"64",x"20",x"C8",x"C1"
		,x"B5",x"EC",x"29",x"01",x"85",x"7F",x"AD",x"02"
		,x"02",x"95",x"B5",x"AD",x"03",x"02",x"95",x"BB"
		,x"A6",x"82",x"A9",x"89",x"95",x"F2",x"AD",x"04"
		,x"02",x"F0",x"10",x"38",x"E9",x"01",x"F0",x"0B"
		,x"D5",x"C7",x"90",x"07",x"A9",x"51",x"8D",x"6C"
		,x"02",x"A9",x"00",x"85",x"D4",x"20",x"0E",x"CE"
		,x"20",x"F8",x"DE",x"50",x"08",x"A9",x"80",x"20"
		,x"97",x"DD",x"4C",x"5E",x"E1",x"20",x"75",x"E2"
		,x"A9",x"80",x"20",x"A6",x"DD",x"F0",x"03",x"4C"
		,x"5E",x"E1",x"4C",x"94",x"C1",x"20",x"9C",x"E2"
		,x"A5",x"D7",x"20",x"C8",x"D4",x"A6",x"82",x"B5"
		,x"C7",x"38",x"E5",x"D4",x"B0",x"03",x"4C",x"02"
		,x"E2",x"18",x"65",x"D7",x"90",x"03",x"69",x"01"
		,x"38",x"20",x"09",x"E0",x"4C",x"38",x"E1",x"A9"
		,x"51",x"20",x"C8",x"C1",x"A5",x"94",x"85",x"89"
		,x"A5",x"95",x"85",x"8A",x"20",x"D0",x"E2",x"D0"
		,x"01",x"60",x"20",x"F1",x"DD",x"20",x"0C",x"DE"
		,x"A5",x"80",x"F0",x"0E",x"20",x"D3",x"E2",x"D0"
		,x"06",x"20",x"1E",x"CF",x"4C",x"DA",x"D2",x"20"
		,x"DA",x"D2",x"A0",x"00",x"B1",x"89",x"85",x"80"
		,x"C8",x"B1",x"89",x"85",x"81",x"4C",x"AF",x"D0"
		,x"20",x"3E",x"DE",x"A0",x"00",x"B1",x"89",x"C5"
		,x"80",x"F0",x"01",x"60",x"C8",x"B1",x"89",x"C5"
		,x"81",x"60",x"20",x"2B",x"DE",x"A0",x"02",x"A9"
		,x"00",x"91",x"94",x"C8",x"D0",x"FB",x"20",x"04"
		,x"E3",x"95",x"C1",x"A8",x"A9",x"FF",x"91",x"94"
		,x"20",x"04",x"E3",x"90",x"F4",x"D0",x"04",x"A9"
		,x"00",x"95",x"C1",x"60",x"A6",x"82",x"B5",x"C1"
		,x"38",x"F0",x"0D",x"18",x"75",x"C7",x"90",x"0B"
		,x"D0",x"06",x"A9",x"02",x"2C",x"CC",x"FE",x"60"
		,x"69",x"01",x"38",x"60",x"20",x"D3",x"D1",x"20"
		,x"CB",x"E1",x"20",x"9C",x"E2",x"20",x"7B",x"CF"
		,x"A5",x"D6",x"85",x"87",x"A5",x"D5",x"85",x"86"
		,x"A9",x"00",x"85",x"88",x"A9",x"00",x"85",x"D4"
		,x"20",x"0E",x"CE",x"20",x"4D",x"EF",x"A4",x"82"
		,x"B6",x"C7",x"CA",x"8A",x"18",x"65",x"D7",x"90"
		,x"0C",x"E6",x"D6",x"E6",x"D6",x"D0",x"06",x"E6"
		,x"D5",x"A9",x"10",x"85",x"D6",x"A5",x"87",x"18"
		,x"69",x"02",x"20",x"E9",x"DE",x"A5",x"D5",x"C9"
		,x"06",x"90",x"05",x"A9",x"52",x"20",x"C8",x"C1"
		,x"A5",x"D6",x"38",x"E5",x"87",x"B0",x"03",x"E9"
		,x"0F",x"18",x"85",x"72",x"A5",x"D5",x"E5",x"86"
		,x"85",x"73",x"A2",x"00",x"86",x"70",x"86",x"71"
		,x"AA",x"20",x"51",x"DF",x"A5",x"71",x"D0",x"07"
		,x"A6",x"70",x"CA",x"D0",x"02",x"E6",x"88",x"CD"
		,x"73",x"02",x"90",x"09",x"D0",x"CD",x"AD",x"72"
		,x"02",x"C5",x"70",x"90",x"C6",x"A9",x"01",x"20"
		,x"F6",x"D4",x"18",x"69",x"01",x"A6",x"82",x"95"
		,x"C1",x"20",x"1E",x"F1",x"20",x"FD",x"DD",x"A5"
		,x"88",x"D0",x"15",x"20",x"5E",x"DE",x"20",x"1E"
		,x"CF",x"20",x"D0",x"D6",x"20",x"1E",x"F1",x"20"
		,x"FD",x"DD",x"20",x"E2",x"E2",x"4C",x"D4",x"E3"
		,x"20",x"1E",x"CF",x"20",x"D0",x"D6",x"20",x"E2"
		,x"E2",x"20",x"19",x"DE",x"20",x"5E",x"DE",x"20"
		,x"0C",x"DE",x"A5",x"80",x"48",x"A5",x"81",x"48"
		,x"20",x"3E",x"DE",x"A5",x"81",x"48",x"A5",x"80"
		,x"48",x"20",x"45",x"DF",x"AA",x"D0",x"0A",x"20"
		,x"4E",x"E4",x"A9",x"10",x"20",x"E9",x"DE",x"E6"
		,x"86",x"68",x"20",x"8D",x"DD",x"68",x"20",x"8D"
		,x"DD",x"68",x"85",x"81",x"68",x"85",x"80",x"F0"
		,x"0F",x"A5",x"86",x"C5",x"D5",x"D0",x"A7",x"20"
		,x"45",x"DF",x"C5",x"D6",x"90",x"A0",x"F0",x"B0"
		,x"20",x"45",x"DF",x"48",x"A9",x"00",x"20",x"DC"
		,x"DE",x"A9",x"00",x"A8",x"91",x"94",x"C8",x"68"
		,x"38",x"E9",x"01",x"91",x"94",x"20",x"6C",x"DE"
		,x"20",x"99",x"D5",x"20",x"F4",x"EE",x"20",x"0E"
		,x"CE",x"20",x"1E",x"CF",x"20",x"F8",x"DE",x"70"
		,x"03",x"4C",x"75",x"E2",x"A9",x"80",x"20",x"97"
		,x"DD",x"A9",x"50",x"20",x"C8",x"C1",x"20",x"1E"
		,x"F1",x"20",x"1E",x"CF",x"20",x"F1",x"DD",x"20"
		,x"93",x"DF",x"48",x"20",x"C1",x"DE",x"A6",x"82"
		,x"B5",x"CD",x"A8",x"68",x"AA",x"A9",x"10",x"20"
		,x"A5",x"DE",x"A9",x"00",x"20",x"DC",x"DE",x"A0"
		,x"02",x"B1",x"94",x"48",x"A9",x"00",x"20",x"C8"
		,x"D4",x"68",x"18",x"69",x"01",x"91",x"94",x"0A"
		,x"69",x"04",x"85",x"89",x"A8",x"38",x"E9",x"02"
		,x"85",x"8A",x"A5",x"80",x"85",x"87",x"91",x"94"
		,x"C8",x"A5",x"81",x"85",x"88",x"91",x"94",x"A0"
		,x"00",x"98",x"91",x"94",x"C8",x"A9",x"11",x"91"
		,x"94",x"A9",x"10",x"20",x"C8",x"D4",x"20",x"50"
		,x"DE",x"20",x"99",x"D5",x"A6",x"82",x"B5",x"CD"
		,x"48",x"20",x"9E",x"DF",x"A6",x"82",x"95",x"CD"
		,x"68",x"AE",x"57",x"02",x"95",x"A7",x"A9",x"00"
		,x"20",x"C8",x"D4",x"A0",x"00",x"A5",x"80",x"91"
		,x"94",x"C8",x"A5",x"81",x"91",x"94",x"4C",x"DE"
		,x"E4",x"20",x"93",x"DF",x"A6",x"82",x"20",x"1B"
		,x"DF",x"A9",x"00",x"20",x"C8",x"D4",x"C6",x"8A"
		,x"C6",x"8A",x"A4",x"89",x"A5",x"87",x"91",x"94"
		,x"C8",x"A5",x"88",x"91",x"94",x"20",x"5E",x"DE"
		,x"20",x"99",x"D5",x"A4",x"8A",x"C0",x"03",x"B0"
		,x"D8",x"4C",x"1E",x"CF",x"00",x"A0",x"4F",x"CB"
		,x"20",x"21",x"22",x"23",x"24",x"27",x"D2",x"45"
		,x"41",x"44",x"89",x"52",x"83",x"20",x"54",x"4F"
		,x"4F",x"20",x"4C",x"41",x"52",x"47",x"C5",x"50"
		,x"8B",x"06",x"20",x"50",x"52",x"45",x"53",x"45"
		,x"4E",x"D4",x"51",x"CF",x"56",x"45",x"52",x"46"
		,x"4C",x"4F",x"57",x"20",x"49",x"4E",x"8B",x"25"
		,x"28",x"8A",x"89",x"26",x"8A",x"20",x"50",x"52"
		,x"4F",x"54",x"45",x"43",x"54",x"20",x"4F",x"CE"
		,x"29",x"88",x"20",x"49",x"44",x"85",x"30",x"31"
		,x"32",x"33",x"34",x"D3",x"59",x"4E",x"54",x"41"
		,x"58",x"89",x"60",x"8A",x"03",x"84",x"63",x"83"
		,x"20",x"45",x"58",x"49",x"53",x"54",x"D3",x"64"
		,x"83",x"20",x"54",x"59",x"50",x"45",x"85",x"65"
		,x"CE",x"4F",x"20",x"42",x"4C",x"4F",x"43",x"CB"
		,x"66",x"67",x"C9",x"4C",x"4C",x"45",x"47",x"41"
		,x"4C",x"20",x"54",x"52",x"41",x"43",x"4B",x"20"
		,x"4F",x"52",x"20",x"53",x"45",x"43",x"54",x"4F"
		,x"D2",x"61",x"83",x"06",x"84",x"39",x"62",x"83"
		,x"06",x"87",x"01",x"83",x"53",x"20",x"53",x"43"
		,x"52",x"41",x"54",x"43",x"48",x"45",x"C4",x"70"
		,x"CE",x"4F",x"20",x"43",x"48",x"41",x"4E",x"4E"
		,x"45",x"CC",x"71",x"C4",x"49",x"52",x"89",x"72"
		,x"88",x"20",x"46",x"55",x"4C",x"CC",x"73",x"C3"
		,x"42",x"4D",x"20",x"44",x"4F",x"53",x"20",x"56"
		,x"32",x"2E",x"36",x"20",x"31",x"35",x"34",x"B1"
		,x"74",x"C4",x"52",x"49",x"56",x"45",x"06",x"20"
		,x"52",x"45",x"41",x"44",x"D9",x"09",x"C5",x"52"
		,x"52",x"4F",x"D2",x"0A",x"D7",x"52",x"49",x"54"
		,x"C5",x"03",x"C6",x"49",x"4C",x"C5",x"04",x"CF"
		,x"50",x"45",x"CE",x"05",x"CD",x"49",x"53",x"4D"
		,x"41",x"54",x"43",x"C8",x"06",x"CE",x"4F",x"D4"
		,x"07",x"C6",x"4F",x"55",x"4E",x"C4",x"08",x"C4"
		,x"49",x"53",x"CB",x"0B",x"D2",x"45",x"43",x"4F"
		,x"52",x"C4",x"48",x"86",x"F9",x"8A",x"0A",x"AA"
		,x"B5",x"06",x"85",x"80",x"B5",x"07",x"85",x"81"
		,x"68",x"29",x"0F",x"F0",x"08",x"C9",x"0F",x"D0"
		,x"06",x"A9",x"74",x"D0",x"08",x"A9",x"06",x"09"
		,x"20",x"AA",x"CA",x"CA",x"8A",x"48",x"AD",x"2A"
		,x"02",x"C9",x"00",x"D0",x"0F",x"A9",x"FF",x"8D"
		,x"2A",x"02",x"68",x"20",x"C7",x"E6",x"20",x"42"
		,x"D0",x"4C",x"48",x"E6",x"68",x"20",x"C7",x"E6"
		,x"20",x"BD",x"C1",x"A9",x"00",x"8D",x"F9",x"02"
		,x"20",x"2C",x"C1",x"20",x"DA",x"D4",x"A9",x"00"
		,x"85",x"A3",x"A2",x"45",x"9A",x"A5",x"84",x"29"
		,x"0F",x"85",x"83",x"C9",x"0F",x"F0",x"31",x"78"
		,x"A5",x"79",x"D0",x"1C",x"A5",x"7A",x"D0",x"10"
		,x"A6",x"83",x"BD",x"2B",x"02",x"C9",x"FF",x"F0"
		,x"1F",x"29",x"0F",x"85",x"82",x"4C",x"8E",x"E6"
		,x"20",x"EB",x"D0",x"EA",x"EA",x"EA",x"D0",x"06"
		,x"20",x"07",x"D1",x"EA",x"EA",x"EA",x"20",x"25"
		,x"D1",x"C9",x"04",x"B0",x"03",x"20",x"27",x"D2"
		,x"4C",x"E7",x"EB",x"AA",x"4C",x"7F",x"C0",x"E0"
		,x"00",x"F0",x"07",x"18",x"69",x"01",x"CA",x"4C"
		,x"9F",x"E6",x"D8",x"AA",x"4A",x"4A",x"4A",x"4A"
		,x"20",x"B4",x"E6",x"8A",x"29",x"0F",x"09",x"30"
		,x"91",x"A5",x"C8",x"60",x"20",x"23",x"C1",x"A9"
		,x"00",x"A0",x"00",x"84",x"80",x"84",x"81",x"A0"
		,x"00",x"A2",x"D5",x"86",x"A5",x"A2",x"02",x"86"
		,x"A6",x"20",x"AB",x"E6",x"A9",x"2C",x"91",x"A5"
		,x"C8",x"AD",x"D5",x"02",x"8D",x"43",x"02",x"8A"
		,x"20",x"06",x"E7",x"A9",x"2C",x"91",x"A5",x"C8"
		,x"A5",x"80",x"20",x"9B",x"E6",x"A9",x"2C",x"91"
		,x"A5",x"C8",x"A5",x"81",x"20",x"9B",x"E6",x"88"
		,x"98",x"18",x"69",x"D5",x"8D",x"49",x"02",x"E6"
		,x"A5",x"A9",x"88",x"85",x"F7",x"60",x"AA",x"A5"
		,x"86",x"48",x"A5",x"87",x"48",x"A9",x"FC",x"85"
		,x"86",x"A9",x"E4",x"85",x"87",x"8A",x"A2",x"00"
		,x"C1",x"86",x"F0",x"21",x"48",x"20",x"75",x"E7"
		,x"90",x"05",x"20",x"75",x"E7",x"90",x"FB",x"A5"
		,x"87",x"C9",x"E6",x"90",x"08",x"D0",x"0A",x"A9"
		,x"0A",x"C5",x"86",x"90",x"04",x"68",x"4C",x"18"
		,x"E7",x"68",x"4C",x"4D",x"E7",x"20",x"67",x"E7"
		,x"90",x"FB",x"20",x"54",x"E7",x"20",x"67",x"E7"
		,x"90",x"F8",x"20",x"54",x"E7",x"68",x"85",x"87"
		,x"68",x"85",x"86",x"60",x"C9",x"20",x"B0",x"0B"
		,x"AA",x"A9",x"20",x"91",x"A5",x"C8",x"8A",x"20"
		,x"06",x"E7",x"60",x"91",x"A5",x"C8",x"60",x"E6"
		,x"86",x"D0",x"02",x"E6",x"87",x"A1",x"86",x"0A"
		,x"A1",x"86",x"29",x"7F",x"60",x"20",x"6D",x"E7"
		,x"E6",x"86",x"D0",x"02",x"E6",x"87",x"60",x"60"
		,x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA"
		,x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA"
		,x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA"
		,x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA",x"EA"
		,x"EA",x"EA",x"60",x"A9",x"8D",x"20",x"68",x"C2"
		,x"20",x"58",x"F2",x"AD",x"78",x"02",x"48",x"A9"
		,x"01",x"8D",x"78",x"02",x"A9",x"FF",x"85",x"86"
		,x"20",x"4F",x"C4",x"AD",x"80",x"02",x"D0",x"05"
		,x"A9",x"39",x"20",x"C8",x"C1",x"68",x"8D",x"78"
		,x"02",x"AD",x"80",x"02",x"85",x"80",x"AD",x"85"
		,x"02",x"85",x"81",x"A9",x"03",x"20",x"77",x"D4"
		,x"A9",x"00",x"85",x"87",x"20",x"39",x"E8",x"85"
		,x"88",x"20",x"4B",x"E8",x"20",x"39",x"E8",x"85"
		,x"89",x"20",x"4B",x"E8",x"A5",x"86",x"F0",x"0A"
		,x"A5",x"88",x"48",x"A5",x"89",x"48",x"A9",x"00"
		,x"85",x"86",x"20",x"39",x"E8",x"85",x"8A",x"20"
		,x"4B",x"E8",x"20",x"39",x"E8",x"A0",x"00",x"91"
		,x"88",x"20",x"4B",x"E8",x"A5",x"88",x"18",x"69"
		,x"01",x"85",x"88",x"90",x"02",x"E6",x"89",x"C6"
		,x"8A",x"D0",x"E7",x"20",x"35",x"CA",x"A5",x"85"
		,x"C5",x"87",x"F0",x"08",x"20",x"3E",x"DE",x"A9"
		,x"50",x"20",x"45",x"E6",x"A5",x"F8",x"D0",x"A8"
		,x"68",x"85",x"89",x"68",x"85",x"88",x"6C",x"88"
		,x"00",x"20",x"35",x"CA",x"A5",x"F8",x"D0",x"08"
		,x"20",x"3E",x"DE",x"A9",x"51",x"20",x"45",x"E6"
		,x"A5",x"85",x"60",x"18",x"65",x"87",x"69",x"00"
		,x"85",x"87",x"60",x"AD",x"01",x"18",x"A9",x"01"
		,x"85",x"7C",x"60",x"78",x"A9",x"00",x"85",x"7C"
		,x"85",x"79",x"85",x"7A",x"A2",x"45",x"9A",x"A9"
		,x"80",x"85",x"F8",x"85",x"7D",x"20",x"B7",x"E9"
		,x"20",x"A5",x"E9",x"AD",x"00",x"18",x"09",x"10"
		,x"8D",x"00",x"18",x"AD",x"00",x"18",x"10",x"57"
		,x"29",x"04",x"D0",x"F7",x"20",x"C9",x"E9",x"C9"
		,x"3F",x"D0",x"06",x"A9",x"00",x"85",x"79",x"F0"
		,x"71",x"C9",x"5F",x"D0",x"06",x"A9",x"00",x"85"
		,x"7A",x"F0",x"67",x"C5",x"78",x"D0",x"0A",x"A9"
		,x"01",x"85",x"7A",x"A9",x"00",x"85",x"79",x"F0"
		,x"29",x"C5",x"77",x"D0",x"0A",x"A9",x"01",x"85"
		,x"79",x"A9",x"00",x"85",x"7A",x"F0",x"1B",x"AA"
		,x"29",x"60",x"C9",x"60",x"D0",x"3F",x"8A",x"85"
		,x"84",x"29",x"0F",x"85",x"83",x"A5",x"84",x"29"
		,x"F0",x"C9",x"E0",x"D0",x"35",x"58",x"20",x"C0"
		,x"DA",x"78",x"2C",x"00",x"18",x"30",x"AD",x"A9"
		,x"00",x"85",x"7D",x"AD",x"00",x"18",x"29",x"EF"
		,x"8D",x"00",x"18",x"A5",x"79",x"F0",x"06",x"20"
		,x"2E",x"EA",x"4C",x"E7",x"EB",x"A5",x"7A",x"F0"
		,x"09",x"20",x"9C",x"E9",x"20",x"AE",x"E9",x"20"
		,x"09",x"E9",x"4C",x"4E",x"EA",x"A9",x"10",x"8D"
		,x"00",x"18",x"2C",x"00",x"18",x"10",x"D0",x"30"
		,x"F9",x"78",x"20",x"EB",x"D0",x"B0",x"06",x"A6"
		,x"82",x"B5",x"F2",x"30",x"01",x"60",x"20",x"59"
		,x"EA",x"20",x"C0",x"E9",x"29",x"01",x"08",x"20"
		,x"B7",x"E9",x"28",x"F0",x"12",x"20",x"59",x"EA"
		,x"20",x"C0",x"E9",x"29",x"01",x"D0",x"F6",x"A6"
		,x"82",x"B5",x"F2",x"29",x"08",x"D0",x"14",x"20"
		,x"59",x"EA",x"20",x"C0",x"E9",x"29",x"01",x"D0"
		,x"F6",x"20",x"59",x"EA",x"20",x"C0",x"E9",x"29"
		,x"01",x"F0",x"F6",x"20",x"AE",x"E9",x"20",x"59"
		,x"EA",x"20",x"C0",x"E9",x"29",x"01",x"D0",x"F3"
		,x"A9",x"08",x"85",x"98",x"20",x"C0",x"E9",x"29"
		,x"01",x"D0",x"36",x"A6",x"82",x"BD",x"3E",x"02"
		,x"6A",x"9D",x"3E",x"02",x"B0",x"05",x"20",x"A5"
		,x"E9",x"D0",x"03",x"20",x"9C",x"E9",x"20",x"B7"
		,x"E9",x"A5",x"23",x"D0",x"03",x"20",x"F3",x"FE"
		,x"20",x"FB",x"FE",x"C6",x"98",x"D0",x"D5",x"20"
		,x"59",x"EA",x"20",x"C0",x"E9",x"29",x"01",x"F0"
		,x"F6",x"58",x"20",x"AA",x"D3",x"78",x"4C",x"0F"
		,x"E9",x"4C",x"4E",x"EA",x"AD",x"00",x"18",x"29"
		,x"FD",x"8D",x"00",x"18",x"60",x"AD",x"00",x"18"
		,x"09",x"02",x"8D",x"00",x"18",x"60",x"AD",x"00"
		,x"18",x"09",x"08",x"8D",x"00",x"18",x"60",x"AD"
		,x"00",x"18",x"29",x"F7",x"8D",x"00",x"18",x"60"
		,x"AD",x"00",x"18",x"CD",x"00",x"18",x"D0",x"F8"
		,x"60",x"A9",x"08",x"85",x"98",x"20",x"59",x"EA"
		,x"20",x"C0",x"E9",x"29",x"04",x"D0",x"F6",x"20"
		,x"9C",x"E9",x"A9",x"01",x"4C",x"20",x"FF",x"20"
		,x"59",x"EA",x"AD",x"0D",x"18",x"29",x"40",x"D0"
		,x"09",x"20",x"C0",x"E9",x"29",x"04",x"F0",x"EF"
		,x"D0",x"19",x"20",x"A5",x"E9",x"A2",x"0A",x"CA"
		,x"D0",x"FD",x"20",x"9C",x"E9",x"20",x"59",x"EA"
		,x"20",x"C0",x"E9",x"29",x"04",x"F0",x"F6",x"A9"
		,x"00",x"85",x"F8",x"AD",x"00",x"18",x"49",x"01"
		,x"4A",x"29",x"02",x"D0",x"F6",x"EA",x"EA",x"EA"
		,x"66",x"85",x"20",x"59",x"EA",x"20",x"C0",x"E9"
		,x"29",x"04",x"F0",x"F6",x"C6",x"98",x"D0",x"E3"
		,x"20",x"A5",x"E9",x"A5",x"85",x"60",x"78",x"20"
		,x"07",x"D1",x"B0",x"05",x"B5",x"F2",x"6A",x"B0"
		,x"0B",x"A5",x"84",x"29",x"F0",x"C9",x"F0",x"F0"
		,x"03",x"4C",x"4E",x"EA",x"20",x"C9",x"E9",x"58"
		,x"20",x"B7",x"CF",x"4C",x"2E",x"EA",x"A9",x"00"
		,x"8D",x"00",x"18",x"4C",x"E7",x"EB",x"4C",x"5B"
		,x"E8",x"A5",x"7D",x"F0",x"06",x"AD",x"00",x"18"
		,x"10",x"09",x"60",x"AD",x"00",x"18",x"10",x"FA"
		,x"4C",x"50",x"FF",x"4C",x"D7",x"E8",x"A2",x"00"
		,x"2C",x"A6",x"6F",x"9A",x"BA",x"A9",x"08",x"0D"
		,x"00",x"1C",x"4C",x"EA",x"FE",x"98",x"18",x"69"
		,x"01",x"D0",x"FC",x"88",x"D0",x"F8",x"AD",x"00"
		,x"1C",x"29",x"F7",x"8D",x"00",x"1C",x"98",x"18"
		,x"69",x"01",x"D0",x"FC",x"88",x"D0",x"F8",x"CA"
		,x"10",x"DB",x"E0",x"FC",x"D0",x"F0",x"F0",x"D4"
		,x"78",x"D8",x"A2",x"FF",x"4C",x"10",x"FF",x"E8"   --EAA0
		,x"A0",x"00",x"A2",x"00",x"8A",x"95",x"00",x"E8"	--EAA8
--		,x"78",x"D8",x"A2",x"FF",x"4C",x"10",x"FF",x"4C"   --EAA0
--		,x"22",x"EB",x"A2",x"00",x"8A",x"95",x"00",x"E8"	--EAA8
		,x"D0",x"FA",x"8A",x"D5",x"00",x"D0",x"B7",x"F6"
		,x"00",x"C8",x"D0",x"FB",x"D5",x"00",x"D0",x"AE"
		,x"94",x"00",x"B5",x"00",x"D0",x"A8",x"E8",x"D0"
		,x"E9",x"E6",x"6F",x"86",x"76",x"A9",x"00",x"85"
		,x"75",x"A8",x"A2",x"20",x"18",x"C6",x"76",x"71"
		,x"75",x"C8",x"D0",x"FB",x"CA",x"D0",x"F6",x"69"
		,x"00",x"AA",x"C5",x"76",x"D0",x"39",x"E0",x"C0"
		,x"D0",x"DF",x"A9",x"01",x"85",x"76",x"E6",x"6F"
		,x"A2",x"07",x"98",x"18",x"65",x"76",x"91",x"75"
		,x"C8",x"D0",x"F7",x"E6",x"76",x"CA",x"D0",x"F2"
		,x"A2",x"07",x"C6",x"76",x"88",x"98",x"18",x"65"
		,x"76",x"D1",x"75",x"D0",x"12",x"49",x"FF",x"91"
		,x"75",x"51",x"75",x"91",x"75",x"D0",x"08",x"98"
		,x"D0",x"EA",x"CA",x"D0",x"E5",x"F0",x"03",x"4C"
		,x"71",x"EA",x"4C",x"49",x"FF",x"AD",x"00",x"1C"
		,x"29",x"F7",x"8D",x"00",x"1C",x"A9",x"01",x"8D"
		,x"0C",x"18",x"A9",x"82",x"8D",x"0D",x"18",x"8D"
		,x"0E",x"18",x"AD",x"00",x"18",x"29",x"60",x"0A"
		,x"2A",x"2A",x"2A",x"09",x"48",x"85",x"78",x"49"
		,x"60",x"85",x"77",x"A2",x"00",x"A0",x"00",x"A9"
		,x"00",x"95",x"99",x"E8",x"B9",x"E0",x"FE",x"95"
		,x"99",x"E8",x"C8",x"C0",x"05",x"D0",x"F0",x"A9"
		,x"00",x"95",x"99",x"E8",x"A9",x"02",x"95",x"99"
		,x"E8",x"A9",x"D5",x"95",x"99",x"E8",x"A9",x"02"
		,x"95",x"99",x"A9",x"FF",x"A2",x"12",x"9D",x"2B"
		,x"02",x"CA",x"10",x"FA",x"A2",x"05",x"95",x"A7"
		,x"95",x"AE",x"95",x"CD",x"CA",x"10",x"F7",x"A9"
		,x"05",x"85",x"AB",x"A9",x"06",x"85",x"AC",x"A9"
		,x"FF",x"85",x"AD",x"85",x"B4",x"A9",x"05",x"8D"
		,x"3B",x"02",x"A9",x"84",x"8D",x"3A",x"02",x"A9"
		,x"0F",x"8D",x"56",x"02",x"A9",x"01",x"85",x"F6"
		,x"A9",x"88",x"85",x"F7",x"A9",x"E0",x"8D",x"4F"
		,x"02",x"A9",x"FF",x"8D",x"50",x"02",x"A9",x"01"
		,x"85",x"1C",x"85",x"1D",x"20",x"63",x"CB",x"20"
		,x"FA",x"CE",x"20",x"59",x"F2",x"A9",x"22",x"85"
		,x"65",x"A9",x"EB",x"85",x"66",x"A9",x"0A",x"85"
		,x"69",x"A9",x"05",x"85",x"6A",x"A9",x"73",x"20"
		,x"C1",x"E6",x"A9",x"00",x"8D",x"00",x"18",x"A9"
		,x"1A",x"8D",x"02",x"18",x"20",x"80",x"E7",x"58"
		,x"AD",x"00",x"18",x"29",x"E5",x"8D",x"00",x"18"
		,x"AD",x"55",x"02",x"F0",x"0A",x"A9",x"00",x"8D"
		,x"55",x"02",x"85",x"67",x"20",x"46",x"C1",x"58"
		,x"A5",x"7C",x"F0",x"03",x"4C",x"50",x"FF",x"58"
		,x"A9",x"0E",x"85",x"72",x"A9",x"00",x"85",x"6F"
		,x"85",x"70",x"A6",x"72",x"BD",x"2B",x"02",x"C9"
		,x"FF",x"F0",x"10",x"29",x"3F",x"85",x"82",x"20"
		,x"93",x"DF",x"AA",x"BD",x"5B",x"02",x"29",x"01"
		,x"AA",x"F6",x"6F",x"C6",x"72",x"10",x"E3",x"A0"
		,x"04",x"B9",x"00",x"00",x"10",x"05",x"29",x"01"
		,x"AA",x"F6",x"6F",x"88",x"10",x"F3",x"78",x"AD"
		,x"00",x"1C",x"29",x"F7",x"48",x"A5",x"7F",x"85"
		,x"86",x"A9",x"00",x"85",x"7F",x"A5",x"6F",x"F0"
		,x"0B",x"A5",x"1C",x"F0",x"03",x"20",x"13",x"D3"
		,x"68",x"09",x"08",x"48",x"E6",x"7F",x"A5",x"70"
		,x"F0",x"0B",x"A5",x"1D",x"F0",x"03",x"20",x"13"
		,x"D3",x"68",x"09",x"00",x"48",x"A5",x"86",x"85"
		,x"7F",x"68",x"AE",x"6C",x"02",x"F0",x"21",x"AD"
		,x"00",x"1C",x"E0",x"80",x"D0",x"03",x"4C",x"8B"
		,x"EC",x"AE",x"05",x"18",x"30",x"12",x"A2",x"A0"
		,x"8E",x"05",x"18",x"CE",x"6C",x"02",x"D0",x"08"
		,x"4D",x"6D",x"02",x"A2",x"10",x"8E",x"6C",x"02"
		,x"8D",x"00",x"1C",x"4C",x"FF",x"EB",x"A9",x"00"
		,x"85",x"83",x"A9",x"01",x"20",x"E2",x"D1",x"A9"
		,x"00",x"20",x"C8",x"D4",x"A6",x"82",x"A9",x"00"
		,x"9D",x"44",x"02",x"20",x"93",x"DF",x"AA",x"A5"
		,x"7F",x"9D",x"5B",x"02",x"A9",x"01",x"20",x"F1"
		,x"CF",x"A9",x"04",x"20",x"F1",x"CF",x"A9",x"01"
		,x"20",x"F1",x"CF",x"20",x"F1",x"CF",x"AD",x"72"
		,x"02",x"20",x"F1",x"CF",x"A9",x"00",x"20",x"F1"
		,x"CF",x"20",x"59",x"ED",x"20",x"93",x"DF",x"0A"
		,x"AA",x"D6",x"99",x"D6",x"99",x"A9",x"00",x"20"
		,x"F1",x"CF",x"A9",x"01",x"20",x"F1",x"CF",x"20"
		,x"F1",x"CF",x"20",x"CE",x"C6",x"90",x"2C",x"AD"
		,x"72",x"02",x"20",x"F1",x"CF",x"AD",x"73",x"02"
		,x"20",x"F1",x"CF",x"20",x"59",x"ED",x"A9",x"00"
		,x"20",x"F1",x"CF",x"D0",x"DD",x"20",x"93",x"DF"
		,x"0A",x"AA",x"A9",x"00",x"95",x"99",x"A9",x"88"
		,x"A4",x"82",x"8D",x"54",x"02",x"99",x"F2",x"00"
		,x"A5",x"85",x"60",x"AD",x"72",x"02",x"20",x"F1"
		,x"CF",x"AD",x"73",x"02",x"20",x"F1",x"CF",x"20"
		,x"59",x"ED",x"20",x"93",x"DF",x"0A",x"AA",x"D6"
		,x"99",x"D6",x"99",x"A9",x"00",x"20",x"F1",x"CF"
		,x"20",x"F1",x"CF",x"20",x"F1",x"CF",x"20",x"93"
		,x"DF",x"0A",x"A8",x"B9",x"99",x"00",x"A6",x"82"
		,x"9D",x"44",x"02",x"DE",x"44",x"02",x"4C",x"0D"
		,x"ED",x"A0",x"00",x"B9",x"B1",x"02",x"20",x"F1"
		,x"CF",x"C8",x"C0",x"1B",x"D0",x"F5",x"60",x"20"
		,x"37",x"D1",x"F0",x"01",x"60",x"85",x"85",x"A4"
		,x"82",x"B9",x"44",x"02",x"F0",x"08",x"A9",x"80"
		,x"99",x"F2",x"00",x"A5",x"85",x"60",x"48",x"20"
		,x"EA",x"EC",x"68",x"60",x"20",x"D1",x"C1",x"20"
		,x"42",x"D0",x"A9",x"40",x"8D",x"F9",x"02",x"20"
		,x"B7",x"EE",x"A9",x"00",x"8D",x"92",x"02",x"20"
		,x"AC",x"C5",x"D0",x"3D",x"A9",x"00",x"85",x"81"
		,x"AD",x"85",x"FE",x"85",x"80",x"20",x"E5",x"ED"
		,x"A9",x"00",x"8D",x"F9",x"02",x"20",x"FF",x"EE"
		,x"4C",x"94",x"C1",x"C8",x"B1",x"94",x"48",x"C8"
		,x"B1",x"94",x"48",x"A0",x"13",x"B1",x"94",x"F0"
		,x"0A",x"85",x"80",x"C8",x"B1",x"94",x"85",x"81"
		,x"20",x"E5",x"ED",x"68",x"85",x"81",x"68",x"85"
		,x"80",x"20",x"E5",x"ED",x"20",x"04",x"C6",x"F0"
		,x"C3",x"A0",x"00",x"B1",x"94",x"30",x"D4",x"20"
		,x"B6",x"C8",x"4C",x"D4",x"ED",x"20",x"5F",x"D5"
		,x"20",x"90",x"EF",x"20",x"75",x"D4",x"A9",x"00"
		,x"20",x"C8",x"D4",x"20",x"37",x"D1",x"85",x"80"
		,x"20",x"37",x"D1",x"85",x"81",x"A5",x"80",x"D0"
		,x"03",x"4C",x"27",x"D2",x"20",x"90",x"EF",x"20"
		,x"4D",x"D4",x"4C",x"EE",x"ED",x"20",x"12",x"C3"
		,x"A5",x"E2",x"10",x"05",x"A9",x"33",x"4C",x"C8"
		,x"C1",x"29",x"01",x"85",x"7F",x"20",x"36",x"FF"
		,x"A5",x"7F",x"0A",x"AA",x"AC",x"7B",x"02",x"CC"
		,x"74",x"02",x"F0",x"1A",x"B9",x"00",x"02",x"95"
		,x"12",x"B9",x"01",x"02",x"95",x"13",x"20",x"07"
		,x"D3",x"A9",x"01",x"85",x"80",x"20",x"2F",x"FF"
		,x"20",x"05",x"F0",x"4C",x"56",x"EE",x"20",x"42"
		,x"D0",x"A6",x"7F",x"BD",x"01",x"01",x"CD",x"D5"
		,x"FE",x"F0",x"03",x"4C",x"72",x"D5",x"20",x"B7"
		,x"EE",x"A5",x"F9",x"A8",x"0A",x"AA",x"AD",x"88"
		,x"FE",x"95",x"99",x"AE",x"7A",x"02",x"A9",x"1B"
		,x"20",x"6E",x"C6",x"A0",x"12",x"A6",x"7F",x"AD"
		,x"D5",x"FE",x"9D",x"01",x"01",x"8A",x"0A",x"AA"
		,x"B5",x"12",x"91",x"94",x"C8",x"B5",x"13",x"91"
		,x"94",x"C8",x"C8",x"A9",x"32",x"91",x"94",x"C8"
		,x"AD",x"D5",x"FE",x"91",x"94",x"A0",x"02",x"91"
		,x"6D",x"AD",x"85",x"FE",x"85",x"80",x"20",x"93"
		,x"EF",x"A9",x"01",x"85",x"81",x"20",x"93",x"EF"
		,x"20",x"FF",x"EE",x"20",x"05",x"F0",x"A0",x"01"
		,x"A9",x"FF",x"91",x"6D",x"20",x"64",x"D4",x"C6"
		,x"81",x"20",x"60",x"D4",x"4C",x"94",x"C1",x"20"
		,x"D1",x"F0",x"A0",x"00",x"A9",x"12",x"91",x"6D"
		,x"C8",x"98",x"91",x"6D",x"C8",x"C8",x"C8",x"A9"
		,x"00",x"85",x"6F",x"85",x"70",x"85",x"71",x"98"
		,x"4A",x"4A",x"20",x"4B",x"F2",x"91",x"6D",x"C8"
		,x"AA",x"38",x"26",x"6F",x"26",x"70",x"26",x"71"
		,x"CA",x"D0",x"F6",x"B5",x"6F",x"91",x"6D",x"C8"
		,x"E8",x"E0",x"03",x"90",x"F6",x"C0",x"90",x"90"
		,x"D6",x"4C",x"75",x"D0",x"20",x"93",x"DF",x"AA"
		,x"BD",x"5B",x"02",x"29",x"01",x"85",x"7F",x"A4"
		,x"7F",x"B9",x"51",x"02",x"D0",x"01",x"60",x"A9"
		,x"00",x"99",x"51",x"02",x"20",x"3A",x"EF",x"A5"
		,x"7F",x"0A",x"48",x"20",x"A5",x"F0",x"68",x"18"
		,x"69",x"01",x"20",x"A5",x"F0",x"A5",x"80",x"48"
		,x"A9",x"01",x"85",x"80",x"0A",x"0A",x"85",x"6D"
		,x"20",x"20",x"F2",x"E6",x"80",x"A5",x"80",x"CD"
		,x"D7",x"FE",x"90",x"F0",x"68",x"85",x"80",x"4C"
		,x"8A",x"D5",x"20",x"0F",x"F1",x"AA",x"20",x"DF"
		,x"F0",x"A6",x"F9",x"BD",x"E0",x"FE",x"85",x"6E"
		,x"A9",x"00",x"85",x"6D",x"60",x"A6",x"7F",x"BD"
		,x"FA",x"02",x"8D",x"72",x"02",x"BD",x"FC",x"02"
		,x"8D",x"73",x"02",x"60",x"20",x"F1",x"EF",x"20"
		,x"CF",x"EF",x"38",x"D0",x"22",x"B1",x"6D",x"1D"
		,x"E9",x"EF",x"91",x"6D",x"20",x"88",x"EF",x"A4"
		,x"6F",x"18",x"B1",x"6D",x"69",x"01",x"91",x"6D"
		,x"A5",x"80",x"CD",x"85",x"FE",x"F0",x"3B",x"FE"
		,x"FA",x"02",x"D0",x"03",x"FE",x"FC",x"02",x"60"
		,x"A6",x"7F",x"A9",x"01",x"9D",x"51",x"02",x"60"
		,x"20",x"F1",x"EF",x"20",x"CF",x"EF",x"F0",x"36"
		,x"B1",x"6D",x"5D",x"E9",x"EF",x"91",x"6D",x"20"
		,x"88",x"EF",x"A4",x"6F",x"B1",x"6D",x"38",x"E9"
		,x"01",x"91",x"6D",x"A5",x"80",x"CD",x"85",x"FE"
		,x"F0",x"0B",x"BD",x"FA",x"02",x"D0",x"03",x"DE"
		,x"FC",x"02",x"DE",x"FA",x"02",x"BD",x"FC",x"02"
		,x"D0",x"0C",x"BD",x"FA",x"02",x"4C",x"93",x"C0"
		,x"EA",x"A9",x"72",x"20",x"C7",x"E6",x"60",x"20"
		,x"11",x"F0",x"98",x"85",x"6F",x"A5",x"81",x"4A"
		,x"4A",x"4A",x"38",x"65",x"6F",x"A8",x"A5",x"81"
		,x"29",x"07",x"AA",x"B1",x"6D",x"3D",x"E9",x"EF"
		,x"60",x"01",x"02",x"04",x"08",x"10",x"20",x"40"
		,x"80",x"A9",x"FF",x"2C",x"F9",x"02",x"F0",x"0C"
		,x"10",x"0A",x"70",x"08",x"A9",x"00",x"8D",x"F9"
		,x"02",x"4C",x"8A",x"D5",x"60",x"20",x"3A",x"EF"
		,x"A0",x"00",x"98",x"91",x"6D",x"C8",x"D0",x"FB"
		,x"60",x"A5",x"6F",x"48",x"A5",x"70",x"48",x"4C"
		,x"5A",x"FF",x"EA",x"F0",x"05",x"A9",x"74",x"20"
		,x"48",x"E6",x"20",x"0F",x"F1",x"85",x"6F",x"8A"
		,x"0A",x"85",x"70",x"AA",x"A5",x"80",x"DD",x"9D"
		,x"02",x"F0",x"0B",x"E8",x"86",x"70",x"DD",x"9D"
		,x"02",x"F0",x"03",x"20",x"5B",x"F0",x"A5",x"70"
		,x"A6",x"7F",x"9D",x"9B",x"02",x"0A",x"0A",x"18"
		,x"69",x"A1",x"85",x"6D",x"A9",x"02",x"69",x"00"
		,x"85",x"6E",x"A0",x"00",x"68",x"85",x"70",x"68"
		,x"85",x"6F",x"60",x"A6",x"6F",x"20",x"DF",x"F0"
		,x"A5",x"7F",x"AA",x"0A",x"1D",x"9B",x"02",x"49"
		,x"01",x"29",x"03",x"85",x"70",x"20",x"A5",x"F0"
		,x"A5",x"F9",x"0A",x"AA",x"A5",x"80",x"0A",x"0A"
		,x"95",x"99",x"A5",x"70",x"0A",x"0A",x"A8",x"A1"
		,x"99",x"99",x"A1",x"02",x"A9",x"00",x"81",x"99"
		,x"F6",x"99",x"C8",x"98",x"29",x"03",x"D0",x"EF"
		,x"A6",x"70",x"A5",x"80",x"9D",x"9D",x"02",x"AD"
		,x"F9",x"02",x"D0",x"03",x"4C",x"8A",x"D5",x"09"
		,x"80",x"8D",x"F9",x"02",x"60",x"A8",x"B9",x"9D"
		,x"02",x"F0",x"25",x"48",x"A9",x"00",x"99",x"9D"
		,x"02",x"A5",x"F9",x"0A",x"AA",x"68",x"0A",x"0A"
		,x"95",x"99",x"98",x"0A",x"0A",x"A8",x"B9",x"A1"
		,x"02",x"81",x"99",x"A9",x"00",x"99",x"A1",x"02"
		,x"F6",x"99",x"C8",x"98",x"29",x"03",x"D0",x"EE"
		,x"60",x"A5",x"7F",x"0A",x"AA",x"A9",x"00",x"9D"
		,x"9D",x"02",x"E8",x"9D",x"9D",x"02",x"60",x"B5"
		,x"A7",x"C9",x"FF",x"D0",x"25",x"8A",x"48",x"20"
		,x"8E",x"D2",x"AA",x"10",x"05",x"A9",x"70",x"20"
		,x"C8",x"C1",x"86",x"F9",x"68",x"A8",x"8A",x"09"
		,x"80",x"99",x"A7",x"00",x"0A",x"AA",x"AD",x"85"
		,x"FE",x"95",x"06",x"A9",x"00",x"95",x"07",x"4C"
		,x"86",x"D5",x"29",x"0F",x"85",x"F9",x"60",x"A9"
		,x"06",x"A6",x"7F",x"D0",x"03",x"18",x"69",x"07"
		,x"60",x"20",x"0F",x"F1",x"AA",x"60",x"20",x"3E"
		,x"DE",x"A9",x"03",x"85",x"6F",x"A9",x"01",x"0D"
		,x"F9",x"02",x"8D",x"F9",x"02",x"A5",x"6F",x"48"
		,x"20",x"11",x"F0",x"68",x"85",x"6F",x"B1",x"6D"
		,x"D0",x"39",x"A5",x"80",x"CD",x"85",x"FE",x"F0"
		,x"19",x"90",x"1C",x"E6",x"80",x"A5",x"80",x"CD"
		,x"D7",x"FE",x"D0",x"E1",x"AE",x"85",x"FE",x"CA"
		,x"86",x"80",x"A9",x"00",x"85",x"81",x"C6",x"6F"
		,x"D0",x"D3",x"A9",x"72",x"20",x"C8",x"C1",x"C6"
		,x"80",x"D0",x"CA",x"AE",x"85",x"FE",x"E8",x"86"
		,x"80",x"A9",x"00",x"85",x"81",x"C6",x"6F",x"D0"
		,x"BC",x"F0",x"E7",x"A5",x"81",x"18",x"65",x"69"
		,x"85",x"81",x"A5",x"80",x"20",x"4B",x"F2",x"8D"
		,x"4E",x"02",x"8D",x"4D",x"02",x"C5",x"81",x"B0"
		,x"0C",x"38",x"A5",x"81",x"ED",x"4E",x"02",x"85"
		,x"81",x"F0",x"02",x"C6",x"81",x"20",x"FA",x"F1"
		,x"F0",x"03",x"4C",x"90",x"EF",x"A9",x"00",x"85"
		,x"81",x"20",x"FA",x"F1",x"D0",x"F4",x"4C",x"F5"
		,x"F1",x"A9",x"01",x"0D",x"F9",x"02",x"8D",x"F9"
		,x"02",x"A5",x"86",x"48",x"A9",x"01",x"85",x"86"
		,x"AD",x"85",x"FE",x"38",x"E5",x"86",x"85",x"80"
		,x"90",x"09",x"F0",x"07",x"20",x"11",x"F0",x"B1"
		,x"6D",x"D0",x"1B",x"AD",x"85",x"FE",x"18",x"65"
		,x"86",x"85",x"80",x"E6",x"86",x"CD",x"D7",x"FE"
		,x"90",x"05",x"A9",x"67",x"20",x"45",x"E6",x"20"
		,x"11",x"F0",x"B1",x"6D",x"F0",x"D2",x"68",x"85"
		,x"86",x"A9",x"00",x"85",x"81",x"20",x"FA",x"F1"
		,x"F0",x"03",x"4C",x"90",x"EF",x"A9",x"71",x"20"
		,x"45",x"E6",x"20",x"11",x"F0",x"98",x"48",x"20"
		,x"20",x"F2",x"A5",x"80",x"20",x"4B",x"F2",x"8D"
		,x"4E",x"02",x"68",x"85",x"6F",x"A5",x"81",x"CD"
		,x"4E",x"02",x"B0",x"09",x"20",x"D5",x"EF",x"D0"
		,x"06",x"E6",x"81",x"D0",x"F0",x"A9",x"00",x"60"
		,x"A5",x"6F",x"48",x"A9",x"00",x"85",x"6F",x"AC"
		,x"86",x"FE",x"88",x"A2",x"07",x"B1",x"6D",x"3D"
		,x"E9",x"EF",x"F0",x"02",x"E6",x"6F",x"CA",x"10"
		,x"F4",x"88",x"D0",x"EF",x"B1",x"6D",x"C5",x"6F"
		,x"D0",x"04",x"68",x"85",x"6F",x"60",x"A9",x"71"
		,x"20",x"45",x"E6",x"AE",x"D6",x"FE",x"DD",x"D6"
		,x"FE",x"CA",x"B0",x"FA",x"BD",x"D1",x"FE",x"60"
		,x"60",x"A9",x"6F",x"8D",x"02",x"1C",x"29",x"F0"
		,x"8D",x"00",x"1C",x"AD",x"0C",x"1C",x"29",x"FE"
		,x"09",x"0E",x"09",x"E0",x"8D",x"0C",x"1C",x"A9"
		,x"41",x"8D",x"0B",x"1C",x"A9",x"00",x"8D",x"06"
		,x"1C",x"A9",x"3A",x"8D",x"07",x"1C",x"8D",x"05"
		,x"1C",x"A9",x"7F",x"8D",x"0E",x"1C",x"A9",x"C0"
		,x"8D",x"0D",x"1C",x"8D",x"0E",x"1C",x"A9",x"FF"
		,x"85",x"3E",x"85",x"51",x"A9",x"08",x"85",x"39"
		,x"A9",x"07",x"85",x"47",x"A9",x"05",x"85",x"62"
		,x"A9",x"FA",x"85",x"63",x"A9",x"C8",x"85",x"64"
		,x"A9",x"04",x"85",x"5E",x"A9",x"04",x"85",x"5F"
		,x"BA",x"86",x"49",x"AD",x"04",x"1C",x"AD",x"0C"
		,x"1C",x"09",x"0E",x"8D",x"0C",x"1C",x"A0",x"05"
		,x"B9",x"00",x"00",x"10",x"2E",x"C9",x"D0",x"D0"
		,x"04",x"98",x"4C",x"70",x"F3",x"29",x"01",x"F0"
		,x"07",x"84",x"3F",x"A9",x"0F",x"4C",x"69",x"F9"
		,x"AA",x"85",x"3D",x"C5",x"3E",x"F0",x"0A",x"20"
		,x"7E",x"F9",x"A5",x"3D",x"85",x"3E",x"4C",x"9C"
		,x"F9",x"A5",x"20",x"30",x"03",x"0A",x"10",x"09"
		,x"4C",x"9C",x"F9",x"88",x"10",x"CA",x"4C",x"9C"
		,x"F9",x"A9",x"20",x"85",x"20",x"A0",x"05",x"84"
		,x"3F",x"20",x"93",x"F3",x"30",x"1A",x"C6",x"3F"
		,x"10",x"F7",x"A4",x"41",x"20",x"95",x"F3",x"A5"
		,x"42",x"85",x"4A",x"06",x"4A",x"A9",x"60",x"85"
		,x"20",x"B1",x"32",x"85",x"22",x"4C",x"9C",x"F9"
		,x"29",x"01",x"C5",x"3D",x"D0",x"E0",x"A5",x"22"
		,x"F0",x"12",x"38",x"F1",x"32",x"F0",x"0D",x"49"
		,x"FF",x"85",x"42",x"E6",x"42",x"A5",x"3F",x"85"
		,x"41",x"4C",x"06",x"F3",x"A2",x"04",x"B1",x"32"
		,x"85",x"40",x"DD",x"D6",x"FE",x"CA",x"B0",x"FA"
		,x"BD",x"D1",x"FE",x"85",x"43",x"8A",x"0A",x"0A"
		,x"0A",x"0A",x"0A",x"85",x"44",x"AD",x"00",x"1C"
		,x"29",x"9F",x"05",x"44",x"8D",x"00",x"1C",x"A6"
		,x"3D",x"A5",x"45",x"C9",x"40",x"F0",x"15",x"C9"
		,x"60",x"F0",x"03",x"4C",x"B1",x"F3",x"A5",x"3F"
		,x"18",x"69",x"03",x"85",x"31",x"A9",x"00",x"85"
		,x"30",x"6C",x"30",x"00",x"A9",x"60",x"85",x"20"
		,x"AD",x"00",x"1C",x"29",x"FC",x"8D",x"00",x"1C"
		,x"A9",x"A4",x"85",x"4A",x"A9",x"01",x"85",x"22"
		,x"4C",x"69",x"F9",x"A4",x"3F",x"B9",x"00",x"00"
		,x"48",x"10",x"10",x"29",x"78",x"85",x"45",x"98"
		,x"0A",x"69",x"06",x"85",x"32",x"98",x"18",x"69"
		,x"03",x"85",x"31",x"A0",x"00",x"84",x"30",x"68"
		,x"60",x"A2",x"5A",x"86",x"4B",x"A2",x"00",x"A9"
		,x"52",x"85",x"24",x"20",x"56",x"F5",x"50",x"FE"
		,x"B8",x"AD",x"01",x"1C",x"C5",x"24",x"D0",x"3F"
		,x"50",x"FE",x"B8",x"AD",x"01",x"1C",x"95",x"25"
		,x"E8",x"E0",x"07",x"D0",x"F3",x"20",x"97",x"F4"
		,x"A0",x"04",x"A9",x"00",x"59",x"16",x"00",x"88"
		,x"10",x"FA",x"C9",x"00",x"D0",x"38",x"A6",x"3E"
		,x"A5",x"18",x"95",x"22",x"A5",x"45",x"C9",x"30"
		,x"F0",x"1E",x"A5",x"3E",x"0A",x"A8",x"B9",x"12"
		,x"00",x"C5",x"16",x"D0",x"1E",x"B9",x"13",x"00"
		,x"C5",x"17",x"D0",x"17",x"4C",x"23",x"F4",x"C6"
		,x"4B",x"D0",x"B0",x"A9",x"02",x"20",x"69",x"F9"
		,x"A5",x"16",x"85",x"12",x"A5",x"17",x"85",x"13"
		,x"A9",x"01",x"2C",x"A9",x"0B",x"2C",x"A9",x"09"
		,x"4C",x"69",x"F9",x"A9",x"7F",x"85",x"4C",x"A5"
		,x"19",x"18",x"69",x"02",x"C5",x"43",x"90",x"02"
		,x"E5",x"43",x"85",x"4D",x"A2",x"05",x"86",x"3F"
		,x"A2",x"FF",x"20",x"93",x"F3",x"10",x"44",x"85"
		,x"44",x"29",x"01",x"C5",x"3E",x"D0",x"3C",x"A0"
		,x"00",x"B1",x"32",x"C5",x"40",x"D0",x"34",x"A5"
		,x"45",x"C9",x"60",x"F0",x"0C",x"A0",x"01",x"38"
		,x"B1",x"32",x"E5",x"4D",x"10",x"03",x"18",x"65"
		,x"43",x"C5",x"4C",x"B0",x"1E",x"48",x"A5",x"45"
		,x"F0",x"14",x"68",x"C9",x"09",x"90",x"14",x"C9"
		,x"0C",x"B0",x"10",x"85",x"4C",x"A5",x"3F",x"AA"
		,x"69",x"03",x"85",x"31",x"D0",x"05",x"68",x"C9"
		,x"06",x"90",x"F0",x"C6",x"3F",x"10",x"B3",x"8A"
		,x"10",x"03",x"4C",x"9C",x"F9",x"86",x"3F",x"20"
		,x"93",x"F3",x"A5",x"45",x"4C",x"CA",x"F4",x"A5"
		,x"30",x"48",x"A5",x"31",x"48",x"A9",x"24",x"85"
		,x"30",x"A9",x"00",x"85",x"31",x"A9",x"00",x"85"
		,x"34",x"20",x"E6",x"F7",x"A5",x"55",x"85",x"18"
		,x"A5",x"54",x"85",x"19",x"A5",x"53",x"85",x"1A"
		,x"20",x"E6",x"F7",x"A5",x"52",x"85",x"17",x"A5"
		,x"53",x"85",x"16",x"68",x"85",x"31",x"68",x"85"
		,x"30",x"60",x"C9",x"00",x"F0",x"03",x"4C",x"6E"
		,x"F5",x"20",x"0A",x"F5",x"50",x"FE",x"B8",x"AD"
		,x"01",x"1C",x"91",x"30",x"C8",x"D0",x"F5",x"A0"
		,x"BA",x"50",x"FE",x"B8",x"AD",x"01",x"1C",x"99"
		,x"00",x"01",x"C8",x"D0",x"F4",x"20",x"E0",x"F8"
		,x"A5",x"38",x"C5",x"47",x"F0",x"05",x"A9",x"04"
		,x"4C",x"69",x"F9",x"20",x"E9",x"F5",x"C5",x"3A"
		,x"F0",x"03",x"A9",x"05",x"2C",x"A9",x"01",x"4C"
		,x"69",x"F9",x"20",x"10",x"F5",x"4C",x"56",x"F5"
		,x"A5",x"3D",x"0A",x"AA",x"B5",x"12",x"85",x"16"
		,x"B5",x"13",x"85",x"17",x"A0",x"00",x"B1",x"32"
		,x"85",x"18",x"C8",x"B1",x"32",x"85",x"19",x"A9"
		,x"00",x"45",x"16",x"45",x"17",x"45",x"18",x"45"
		,x"19",x"85",x"1A",x"20",x"34",x"F9",x"A2",x"5A"
		,x"20",x"56",x"F5",x"A0",x"00",x"50",x"FE",x"B8"
		,x"AD",x"01",x"1C",x"D9",x"24",x"00",x"D0",x"06"
		,x"C8",x"C0",x"08",x"D0",x"F0",x"60",x"CA",x"D0"
		,x"E7",x"A9",x"02",x"4C",x"69",x"F9",x"A9",x"D0"
		,x"8D",x"05",x"18",x"A9",x"03",x"2C",x"05",x"18"
		,x"10",x"F1",x"2C",x"00",x"1C",x"30",x"F6",x"AD"
		,x"01",x"1C",x"B8",x"A0",x"00",x"60",x"C9",x"10"
		,x"F0",x"03",x"4C",x"91",x"F6",x"20",x"E9",x"F5"
		,x"85",x"3A",x"AD",x"00",x"1C",x"29",x"10",x"D0"
		,x"05",x"A9",x"08",x"4C",x"69",x"F9",x"20",x"8F"
		,x"F7",x"20",x"10",x"F5",x"A2",x"09",x"50",x"FE"
		,x"B8",x"CA",x"D0",x"FA",x"A9",x"FF",x"8D",x"03"
		,x"1C",x"AD",x"0C",x"1C",x"29",x"1F",x"09",x"C0"
		,x"8D",x"0C",x"1C",x"A9",x"FF",x"A2",x"05",x"8D"
		,x"01",x"1C",x"B8",x"50",x"FE",x"B8",x"CA",x"D0"
		,x"FA",x"A0",x"BB",x"B9",x"00",x"01",x"50",x"FE"
		,x"B8",x"8D",x"01",x"1C",x"C8",x"D0",x"F4",x"B1"
		,x"30",x"50",x"FE",x"B8",x"8D",x"01",x"1C",x"C8"
		,x"D0",x"F5",x"50",x"FE",x"AD",x"0C",x"1C",x"09"
		,x"E0",x"8D",x"0C",x"1C",x"A9",x"00",x"8D",x"03"
		,x"1C",x"20",x"F2",x"F5",x"A4",x"3F",x"B9",x"00"
		,x"00",x"49",x"30",x"99",x"00",x"00",x"4C",x"B1"
		,x"F3",x"A9",x"00",x"A8",x"51",x"30",x"C8",x"D0"
		,x"FB",x"60",x"A9",x"00",x"85",x"2E",x"85",x"30"
		,x"85",x"4F",x"A5",x"31",x"85",x"4E",x"A9",x"01"
		,x"85",x"31",x"85",x"2F",x"A9",x"BB",x"85",x"34"
		,x"85",x"36",x"20",x"E6",x"F7",x"A5",x"52",x"85"
		,x"38",x"A4",x"36",x"A5",x"53",x"91",x"2E",x"C8"
		,x"A5",x"54",x"91",x"2E",x"C8",x"A5",x"55",x"91"
		,x"2E",x"C8",x"84",x"36",x"20",x"E6",x"F7",x"A4"
		,x"36",x"A5",x"52",x"91",x"2E",x"C8",x"A5",x"53"
		,x"91",x"2E",x"C8",x"F0",x"0E",x"A5",x"54",x"91"
		,x"2E",x"C8",x"A5",x"55",x"91",x"2E",x"C8",x"84"
		,x"36",x"D0",x"E1",x"A5",x"54",x"91",x"30",x"C8"
		,x"A5",x"55",x"91",x"30",x"C8",x"84",x"36",x"20"
		,x"E6",x"F7",x"A4",x"36",x"A5",x"52",x"91",x"30"
		,x"C8",x"A5",x"53",x"91",x"30",x"C8",x"A5",x"54"
		,x"91",x"30",x"C8",x"A5",x"55",x"91",x"30",x"C8"
		,x"84",x"36",x"C0",x"BB",x"90",x"E1",x"A9",x"45"
		,x"85",x"2E",x"A5",x"31",x"85",x"2F",x"A0",x"BA"
		,x"B1",x"30",x"91",x"2E",x"88",x"D0",x"F9",x"B1"
		,x"30",x"91",x"2E",x"A2",x"BB",x"BD",x"00",x"01"
		,x"91",x"30",x"C8",x"E8",x"D0",x"F7",x"86",x"50"
		,x"60",x"C9",x"20",x"F0",x"03",x"4C",x"CA",x"F6"
		,x"20",x"E9",x"F5",x"85",x"3A",x"20",x"8F",x"F7"
		,x"20",x"0A",x"F5",x"A0",x"BB",x"B9",x"00",x"01"
		,x"50",x"FE",x"B8",x"4D",x"01",x"1C",x"D0",x"15"
		,x"C8",x"D0",x"F2",x"B1",x"30",x"50",x"FE",x"B8"
		,x"4D",x"01",x"1C",x"D0",x"08",x"C8",x"C0",x"FD"
		,x"D0",x"F1",x"4C",x"18",x"F4",x"A9",x"07",x"4C"
		,x"69",x"F9",x"20",x"10",x"F5",x"4C",x"18",x"F4"
		,x"A9",x"00",x"85",x"57",x"85",x"5A",x"A4",x"34"
		,x"A5",x"52",x"29",x"F0",x"4A",x"4A",x"4A",x"4A"
		,x"AA",x"BD",x"7F",x"F7",x"0A",x"0A",x"0A",x"85"
		,x"56",x"A5",x"52",x"29",x"0F",x"AA",x"BD",x"7F"
		,x"F7",x"6A",x"66",x"57",x"6A",x"66",x"57",x"29"
		,x"07",x"05",x"56",x"91",x"30",x"C8",x"A5",x"53"
		,x"29",x"F0",x"4A",x"4A",x"4A",x"4A",x"AA",x"BD"
		,x"7F",x"F7",x"0A",x"05",x"57",x"85",x"57",x"A5"
		,x"53",x"29",x"0F",x"AA",x"BD",x"7F",x"F7",x"2A"
		,x"2A",x"2A",x"2A",x"85",x"58",x"2A",x"29",x"01"
		,x"05",x"57",x"91",x"30",x"C8",x"A5",x"54",x"29"
		,x"F0",x"4A",x"4A",x"4A",x"4A",x"AA",x"BD",x"7F"
		,x"F7",x"18",x"6A",x"05",x"58",x"91",x"30",x"C8"
		,x"6A",x"29",x"80",x"85",x"59",x"A5",x"54",x"29"
		,x"0F",x"AA",x"BD",x"7F",x"F7",x"0A",x"0A",x"29"
		,x"7C",x"05",x"59",x"85",x"59",x"A5",x"55",x"29"
		,x"F0",x"4A",x"4A",x"4A",x"4A",x"AA",x"BD",x"7F"
		,x"F7",x"6A",x"66",x"5A",x"6A",x"66",x"5A",x"6A"
		,x"66",x"5A",x"29",x"03",x"05",x"59",x"91",x"30"
		,x"C8",x"D0",x"04",x"A5",x"2F",x"85",x"31",x"A5"
		,x"55",x"29",x"0F",x"AA",x"BD",x"7F",x"F7",x"05"
		,x"5A",x"91",x"30",x"C8",x"84",x"34",x"60",x"0A"
		,x"0B",x"12",x"13",x"0E",x"0F",x"16",x"17",x"09"
		,x"19",x"1A",x"1B",x"0D",x"1D",x"1E",x"15",x"A9"
		,x"00",x"85",x"30",x"85",x"2E",x"85",x"36",x"A9"
		,x"BB",x"85",x"34",x"85",x"50",x"A5",x"31",x"85"
		,x"2F",x"A9",x"01",x"85",x"31",x"A5",x"47",x"85"
		,x"52",x"A4",x"36",x"B1",x"2E",x"85",x"53",x"C8"
		,x"B1",x"2E",x"85",x"54",x"C8",x"B1",x"2E",x"85"
		,x"55",x"C8",x"84",x"36",x"20",x"D0",x"F6",x"A4"
		,x"36",x"B1",x"2E",x"85",x"52",x"C8",x"F0",x"11"
		,x"B1",x"2E",x"85",x"53",x"C8",x"B1",x"2E",x"85"
		,x"54",x"C8",x"B1",x"2E",x"85",x"55",x"C8",x"D0"
		,x"E1",x"A5",x"3A",x"85",x"53",x"A9",x"00",x"85"
		,x"54",x"85",x"55",x"4C",x"D0",x"F6",x"A4",x"34"
		,x"B1",x"30",x"29",x"F8",x"4A",x"4A",x"4A",x"85"
		,x"56",x"B1",x"30",x"29",x"07",x"0A",x"0A",x"85"
		,x"57",x"C8",x"D0",x"06",x"A5",x"4E",x"85",x"31"
		,x"A4",x"4F",x"B1",x"30",x"29",x"C0",x"2A",x"2A"
		,x"2A",x"05",x"57",x"85",x"57",x"B1",x"30",x"29"
		,x"3E",x"4A",x"85",x"58",x"B1",x"30",x"29",x"01"
		,x"0A",x"0A",x"0A",x"0A",x"85",x"59",x"C8",x"B1"
		,x"30",x"29",x"F0",x"4A",x"4A",x"4A",x"4A",x"05"
		,x"59",x"85",x"59",x"B1",x"30",x"29",x"0F",x"0A"
		,x"85",x"5A",x"C8",x"B1",x"30",x"29",x"80",x"18"
		,x"2A",x"2A",x"29",x"01",x"05",x"5A",x"85",x"5A"
		,x"B1",x"30",x"29",x"7C",x"4A",x"4A",x"85",x"5B"
		,x"B1",x"30",x"29",x"03",x"0A",x"0A",x"0A",x"85"
		,x"5C",x"C8",x"D0",x"06",x"A5",x"4E",x"85",x"31"
		,x"A4",x"4F",x"B1",x"30",x"29",x"E0",x"2A",x"2A"
		,x"2A",x"2A",x"05",x"5C",x"85",x"5C",x"B1",x"30"
		,x"29",x"1F",x"85",x"5D",x"C8",x"84",x"34",x"A6"
		,x"56",x"BD",x"A0",x"F8",x"A6",x"57",x"1D",x"C0"
		,x"F8",x"85",x"52",x"A6",x"58",x"BD",x"A0",x"F8"
		,x"A6",x"59",x"1D",x"C0",x"F8",x"85",x"53",x"A6"
		,x"5A",x"BD",x"A0",x"F8",x"A6",x"5B",x"1D",x"C0"
		,x"F8",x"85",x"54",x"A6",x"5C",x"BD",x"A0",x"F8"
		,x"A6",x"5D",x"1D",x"C0",x"F8",x"85",x"55",x"60"
		,x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"
		,x"FF",x"80",x"00",x"10",x"FF",x"C0",x"40",x"50"
		,x"FF",x"FF",x"20",x"30",x"FF",x"F0",x"60",x"70"
		,x"FF",x"90",x"A0",x"B0",x"FF",x"D0",x"E0",x"FF"
		,x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF"
		,x"FF",x"08",x"00",x"01",x"FF",x"0C",x"04",x"05"
		,x"FF",x"FF",x"02",x"03",x"FF",x"0F",x"06",x"07"
		,x"FF",x"09",x"0A",x"0B",x"FF",x"0D",x"0E",x"FF"
		,x"A9",x"00",x"85",x"34",x"85",x"2E",x"85",x"36"
		,x"A9",x"01",x"85",x"4E",x"A9",x"BA",x"85",x"4F"
		,x"A5",x"31",x"85",x"2F",x"20",x"E6",x"F7",x"A5"
		,x"52",x"85",x"38",x"A4",x"36",x"A5",x"53",x"91"
		,x"2E",x"C8",x"A5",x"54",x"91",x"2E",x"C8",x"A5"
		,x"55",x"91",x"2E",x"C8",x"84",x"36",x"20",x"E6"
		,x"F7",x"A4",x"36",x"A5",x"52",x"91",x"2E",x"C8"
		,x"F0",x"11",x"A5",x"53",x"91",x"2E",x"C8",x"A5"
		,x"54",x"91",x"2E",x"C8",x"A5",x"55",x"91",x"2E"
		,x"C8",x"D0",x"E1",x"A5",x"53",x"85",x"3A",x"A5"
		,x"2F",x"85",x"31",x"60",x"A5",x"31",x"85",x"2F"
		,x"A9",x"00",x"85",x"31",x"A9",x"24",x"85",x"34"
		,x"A5",x"39",x"85",x"52",x"A5",x"1A",x"85",x"53"
		,x"A5",x"19",x"85",x"54",x"A5",x"18",x"85",x"55"
		,x"20",x"D0",x"F6",x"A5",x"17",x"85",x"52",x"A5"
		,x"16",x"85",x"53",x"A9",x"00",x"85",x"54",x"85"
		,x"55",x"20",x"D0",x"F6",x"A5",x"2F",x"85",x"31"
		,x"60",x"A4",x"3F",x"99",x"00",x"00",x"A5",x"50"
		,x"F0",x"03",x"20",x"F2",x"F5",x"20",x"8F",x"F9"
		,x"A6",x"49",x"9A",x"4C",x"BE",x"F2",x"A9",x"A0"
		,x"85",x"20",x"AD",x"00",x"1C",x"09",x"04",x"8D"
		,x"00",x"1C",x"A9",x"3C",x"85",x"48",x"60",x"A6"
		,x"3E",x"A5",x"20",x"09",x"10",x"85",x"20",x"A9"
		,x"FF",x"85",x"48",x"60",x"AD",x"07",x"1C",x"8D"
		,x"05",x"1C",x"AD",x"00",x"1C",x"29",x"10",x"C5"
		,x"1E",x"85",x"1E",x"F0",x"04",x"A9",x"01",x"85"
		,x"1C",x"AD",x"FE",x"02",x"F0",x"15",x"C9",x"02"
		,x"D0",x"07",x"A9",x"00",x"8D",x"FE",x"02",x"F0"
		,x"0A",x"85",x"4A",x"A9",x"02",x"8D",x"FE",x"02"
		,x"4C",x"2E",x"FA",x"A6",x"3E",x"30",x"07",x"A5"
		,x"20",x"A8",x"C9",x"20",x"D0",x"03",x"4C",x"BE"
		,x"FA",x"C6",x"48",x"D0",x"1D",x"98",x"10",x"04"
		,x"29",x"7F",x"85",x"20",x"29",x"10",x"F0",x"12"
		,x"AD",x"00",x"1C",x"29",x"FB",x"8D",x"00",x"1C"
		,x"A9",x"FF",x"85",x"3E",x"A9",x"00",x"85",x"20"
		,x"F0",x"DC",x"98",x"29",x"40",x"D0",x"03",x"4C"
		,x"BE",x"FA",x"6C",x"62",x"00",x"A5",x"4A",x"10"
		,x"05",x"49",x"FF",x"18",x"69",x"01",x"C5",x"64"
		,x"B0",x"0A",x"A9",x"3B",x"85",x"62",x"A9",x"FA"
		,x"85",x"63",x"D0",x"12",x"E5",x"5E",x"E5",x"5E"
		,x"85",x"61",x"A5",x"5E",x"85",x"60",x"A9",x"7B"
		,x"85",x"62",x"A9",x"FA",x"85",x"63",x"A5",x"4A"
		,x"10",x"31",x"E6",x"4A",x"AE",x"00",x"1C",x"CA"
		,x"4C",x"69",x"FA",x"A5",x"4A",x"D0",x"EF",x"A9"
		,x"4E",x"85",x"62",x"A9",x"FA",x"85",x"63",x"A9"
		,x"05",x"85",x"60",x"4C",x"BE",x"FA",x"C6",x"60"
		,x"D0",x"6C",x"A5",x"20",x"29",x"BF",x"85",x"20"
		,x"A9",x"05",x"85",x"62",x"A9",x"FA",x"85",x"63"
		,x"4C",x"BE",x"FA",x"C6",x"4A",x"AE",x"00",x"1C"
		,x"E8",x"8A",x"29",x"03",x"85",x"4B",x"AD",x"00"
		,x"1C",x"29",x"FC",x"05",x"4B",x"8D",x"00",x"1C"
		,x"4C",x"BE",x"FA",x"38",x"AD",x"07",x"1C",x"E5"
		,x"5F",x"8D",x"05",x"1C",x"C6",x"60",x"D0",x"0C"
		,x"A5",x"5E",x"85",x"60",x"A9",x"97",x"85",x"62"
		,x"A9",x"FA",x"85",x"63",x"4C",x"2E",x"FA",x"C6"
		,x"61",x"D0",x"F9",x"A9",x"A5",x"85",x"62",x"A9"
		,x"FA",x"85",x"63",x"D0",x"EF",x"AD",x"07",x"1C"
		,x"18",x"65",x"5F",x"8D",x"05",x"1C",x"C6",x"60"
		,x"D0",x"E2",x"A9",x"4E",x"85",x"62",x"A9",x"FA"
		,x"85",x"63",x"A9",x"05",x"85",x"60",x"AD",x"0C"
		,x"1C",x"29",x"FD",x"8D",x"0C",x"1C",x"60",x"A5"
		,x"51",x"10",x"2A",x"A6",x"3D",x"A9",x"60",x"95"
		,x"20",x"A9",x"01",x"95",x"22",x"85",x"51",x"A9"
		,x"A4",x"85",x"4A",x"AD",x"00",x"1C",x"29",x"FC"
		,x"8D",x"00",x"1C",x"A9",x"0A",x"8D",x"20",x"06"
		,x"A9",x"A0",x"8D",x"21",x"06",x"A9",x"0F",x"8D"
		,x"22",x"06",x"4C",x"9C",x"F9",x"A0",x"00",x"D1"
		,x"32",x"F0",x"05",x"91",x"32",x"4C",x"9C",x"F9"
		,x"AD",x"00",x"1C",x"29",x"10",x"D0",x"05",x"A9"
		,x"08",x"4C",x"D3",x"FD",x"20",x"A3",x"FD",x"20"
		,x"C3",x"FD",x"A9",x"55",x"8D",x"01",x"1C",x"20"
		,x"C3",x"FD",x"20",x"00",x"FE",x"20",x"56",x"F5"
		,x"A9",x"40",x"0D",x"0B",x"18",x"8D",x"0B",x"18"
		,x"A9",x"62",x"8D",x"06",x"18",x"A9",x"00",x"8D"
		,x"07",x"18",x"8D",x"05",x"18",x"A0",x"00",x"A2"
		,x"00",x"2C",x"00",x"1C",x"30",x"FB",x"2C",x"00"
		,x"1C",x"10",x"FB",x"AD",x"04",x"18",x"2C",x"00"
		,x"1C",x"10",x"11",x"AD",x"0D",x"18",x"0A",x"10"
		,x"F5",x"E8",x"D0",x"EF",x"C8",x"D0",x"EC",x"A9"
		,x"02",x"4C",x"D3",x"FD",x"86",x"71",x"84",x"72"
		,x"A2",x"00",x"A0",x"00",x"AD",x"04",x"18",x"2C"
		,x"00",x"1C",x"30",x"11",x"AD",x"0D",x"18",x"0A"
		,x"10",x"F5",x"E8",x"D0",x"EF",x"C8",x"D0",x"EC"
		,x"A9",x"02",x"4C",x"D3",x"FD",x"38",x"8A",x"E5"
		,x"71",x"AA",x"85",x"70",x"98",x"E5",x"72",x"A8"
		,x"85",x"71",x"10",x"0B",x"49",x"FF",x"A8",x"8A"
		,x"49",x"FF",x"AA",x"E8",x"D0",x"01",x"C8",x"98"
		,x"D0",x"04",x"E0",x"04",x"90",x"18",x"06",x"70"
		,x"26",x"71",x"18",x"A5",x"70",x"6D",x"21",x"06"
		,x"8D",x"21",x"06",x"A5",x"71",x"6D",x"22",x"06"
		,x"8D",x"22",x"06",x"4C",x"0C",x"FB",x"A2",x"00"
		,x"A0",x"00",x"B8",x"AD",x"00",x"1C",x"10",x"0E"
		,x"50",x"F9",x"B8",x"E8",x"D0",x"F5",x"C8",x"D0"
		,x"F2",x"A9",x"03",x"4C",x"D3",x"FD",x"8A",x"0A"
		,x"8D",x"25",x"06",x"98",x"2A",x"8D",x"24",x"06"
		,x"A9",x"BF",x"2D",x"0B",x"18",x"8D",x"0B",x"18"
		,x"A9",x"66",x"8D",x"26",x"06",x"A6",x"43",x"A0"
		,x"00",x"98",x"18",x"6D",x"26",x"06",x"90",x"01"
		,x"C8",x"C8",x"CA",x"D0",x"F5",x"49",x"FF",x"38"
		,x"69",x"00",x"18",x"6D",x"25",x"06",x"B0",x"03"
		,x"CE",x"24",x"06",x"AA",x"98",x"49",x"FF",x"38"
		,x"69",x"00",x"18",x"6D",x"24",x"06",x"10",x"05"
		,x"A9",x"04",x"4C",x"D3",x"FD",x"A8",x"8A",x"A2"
		,x"00",x"38",x"E5",x"43",x"B0",x"03",x"88",x"30"
		,x"03",x"E8",x"D0",x"F5",x"8E",x"26",x"06",x"E0"
		,x"04",x"B0",x"05",x"A9",x"05",x"4C",x"D3",x"FD"
		,x"18",x"65",x"43",x"8D",x"27",x"06",x"A9",x"00"
		,x"8D",x"28",x"06",x"A0",x"00",x"A6",x"3D",x"A5"
		,x"39",x"99",x"00",x"03",x"C8",x"C8",x"AD",x"28"
		,x"06",x"99",x"00",x"03",x"C8",x"A5",x"51",x"99"
		,x"00",x"03",x"C8",x"B5",x"13",x"99",x"00",x"03"
		,x"C8",x"B5",x"12",x"99",x"00",x"03",x"C8",x"A9"
		,x"0F",x"99",x"00",x"03",x"C8",x"99",x"00",x"03"
		,x"C8",x"A9",x"00",x"59",x"FA",x"02",x"59",x"FB"
		,x"02",x"59",x"FC",x"02",x"59",x"FD",x"02",x"99"
		,x"F9",x"02",x"EE",x"28",x"06",x"AD",x"28",x"06"
		,x"C5",x"43",x"90",x"BB",x"98",x"48",x"E8",x"8A"
		,x"9D",x"00",x"05",x"E8",x"D0",x"FA",x"A9",x"03"
		,x"85",x"31",x"20",x"30",x"FE",x"68",x"A8",x"88"
		,x"20",x"E5",x"FD",x"20",x"F5",x"FD",x"A9",x"05"
		,x"85",x"31",x"20",x"E9",x"F5",x"85",x"3A",x"20"
		,x"8F",x"F7",x"A9",x"00",x"85",x"32",x"20",x"4E"
		,x"C0",x"A9",x"FF",x"8D",x"01",x"1C",x"A2",x"05"
		,x"50",x"FE",x"B8",x"CA",x"D0",x"FA",x"A2",x"0A"
		,x"A4",x"32",x"50",x"FE",x"B8",x"B9",x"00",x"03"
		,x"8D",x"01",x"1C",x"C8",x"CA",x"D0",x"F3",x"A2"
		,x"09",x"50",x"FE",x"B8",x"A9",x"55",x"8D",x"01"
		,x"1C",x"CA",x"D0",x"F5",x"A9",x"FF",x"A2",x"05"
		,x"50",x"FE",x"B8",x"8D",x"01",x"1C",x"CA",x"D0"
		,x"F7",x"A2",x"BB",x"50",x"FE",x"B8",x"BD",x"00"
		,x"01",x"8D",x"01",x"1C",x"E8",x"D0",x"F4",x"A0"
		,x"00",x"50",x"FE",x"B8",x"B1",x"30",x"8D",x"01"
		,x"1C",x"C8",x"D0",x"F5",x"A9",x"55",x"AE",x"26"
		,x"06",x"50",x"FE",x"B8",x"8D",x"01",x"1C",x"CA"
		,x"D0",x"F7",x"A5",x"32",x"18",x"69",x"0A",x"85"
		,x"32",x"CE",x"28",x"06",x"D0",x"93",x"50",x"FE"
		,x"B8",x"50",x"FE",x"B8",x"20",x"00",x"FE",x"A9"
		,x"C8",x"8D",x"23",x"06",x"A9",x"00",x"85",x"30"
		,x"A9",x"03",x"85",x"31",x"A5",x"43",x"8D",x"28"
		,x"06",x"20",x"56",x"F5",x"A2",x"0A",x"A0",x"00"
		,x"50",x"FE",x"B8",x"AD",x"01",x"1C",x"D1",x"30"
		,x"D0",x"0E",x"C8",x"CA",x"D0",x"F2",x"18",x"A5"
		,x"30",x"69",x"0A",x"85",x"30",x"4C",x"62",x"FD"
		,x"CE",x"23",x"06",x"D0",x"CF",x"A9",x"06",x"4C"
		,x"D3",x"FD",x"20",x"56",x"F5",x"A0",x"BB",x"50"
		,x"FE",x"B8",x"AD",x"01",x"1C",x"D9",x"00",x"01"
		,x"D0",x"E6",x"C8",x"D0",x"F2",x"A2",x"FC",x"50"
		,x"FE",x"B8",x"AD",x"01",x"1C",x"D9",x"00",x"05"
		,x"D0",x"D6",x"C8",x"CA",x"D0",x"F1",x"CE",x"28"
		,x"06",x"D0",x"AE",x"E6",x"51",x"A5",x"51",x"C9"
		,x"24",x"B0",x"03",x"4C",x"9C",x"F9",x"A9",x"FF"
		,x"85",x"51",x"A9",x"00",x"85",x"50",x"A9",x"01"
		,x"4C",x"69",x"F9",x"AD",x"0C",x"1C",x"29",x"1F"
		,x"09",x"C0",x"8D",x"0C",x"1C",x"A9",x"FF",x"8D"
		,x"03",x"1C",x"8D",x"01",x"1C",x"A2",x"28",x"A0"
		,x"00",x"50",x"FE",x"B8",x"88",x"D0",x"FA",x"CA"
		,x"D0",x"F7",x"60",x"AE",x"21",x"06",x"AC",x"22"
		,x"06",x"50",x"FE",x"B8",x"CA",x"D0",x"FA",x"88"
		,x"10",x"F7",x"60",x"CE",x"20",x"06",x"F0",x"03"
		,x"4C",x"9C",x"F9",x"A0",x"FF",x"84",x"51",x"C8"
		,x"84",x"50",x"4C",x"69",x"F9",x"B9",x"00",x"03"
		,x"99",x"45",x"03",x"88",x"D0",x"F7",x"AD",x"00"
		,x"03",x"8D",x"45",x"03",x"60",x"A0",x"44",x"B9"
		,x"BB",x"01",x"91",x"30",x"88",x"10",x"F8",x"60"
		,x"AD",x"0C",x"1C",x"09",x"E0",x"8D",x"0C",x"1C"
		,x"A9",x"00",x"8D",x"03",x"1C",x"60",x"AD",x"0C"
		,x"1C",x"29",x"1F",x"09",x"C0",x"8D",x"0C",x"1C"
		,x"A9",x"FF",x"8D",x"03",x"1C",x"A9",x"55",x"8D"
		,x"01",x"1C",x"A2",x"28",x"A0",x"00",x"50",x"FE"
		,x"B8",x"88",x"D0",x"FA",x"CA",x"D0",x"F7",x"60"
		,x"A9",x"00",x"85",x"30",x"85",x"2E",x"85",x"36"
		,x"A9",x"BB",x"85",x"34",x"A5",x"31",x"85",x"2F"
		,x"A9",x"01",x"85",x"31",x"A4",x"36",x"B1",x"2E"
		,x"85",x"52",x"C8",x"B1",x"2E",x"85",x"53",x"C8"
		,x"B1",x"2E",x"85",x"54",x"C8",x"B1",x"2E",x"85"
		,x"55",x"C8",x"F0",x"08",x"84",x"36",x"20",x"D0"
		,x"F6",x"4C",x"44",x"FE",x"4C",x"D0",x"F6",x"48"
		,x"8A",x"48",x"98",x"48",x"AD",x"0D",x"18",x"29"
		,x"02",x"F0",x"03",x"20",x"53",x"E8",x"AD",x"0D"
		,x"1C",x"0A",x"10",x"03",x"20",x"B0",x"F2",x"68"
		,x"A8",x"68",x"AA",x"68",x"40",x"12",x"04",x"04"
		,x"90",x"56",x"49",x"44",x"4D",x"42",x"55",x"50"
		,x"26",x"43",x"52",x"53",x"4E",x"84",x"05",x"C1"
		,x"F8",x"1B",x"5C",x"07",x"A3",x"F0",x"88",x"23"
		,x"0D",x"ED",x"D0",x"C8",x"CA",x"CC",x"CB",x"E2"
		,x"E7",x"C8",x"CA",x"C8",x"EE",x"51",x"DD",x"1C"
		,x"9E",x"1C",x"52",x"57",x"41",x"4D",x"44",x"53"
		,x"50",x"55",x"4C",x"44",x"53",x"50",x"55",x"52"
		,x"45",x"45",x"52",x"53",x"45",x"4C",x"51",x"47"
		,x"52",x"4C",x"08",x"00",x"00",x"3F",x"7F",x"BF"
		,x"FF",x"11",x"12",x"13",x"15",x"41",x"04",x"24"
		,x"1F",x"19",x"12",x"01",x"FF",x"FF",x"01",x"00"
		,x"03",x"04",x"05",x"06",x"07",x"07",x"79",x"6C"
		,x"65",x"00",x"8D",x"00",x"1C",x"8D",x"02",x"1C"
		,x"4C",x"7D",x"EA",x"8A",x"A2",x"05",x"CA",x"D0"
		,x"FD",x"AA",x"60",x"20",x"AE",x"E9",x"4C",x"9C"
		,x"E9",x"AD",x"02",x"02",x"C9",x"2D",x"F0",x"05"
		,x"38",x"E9",x"2B",x"D0",x"DA",x"85",x"23",x"60"
		,x"8E",x"03",x"18",x"A9",x"02",x"8D",x"00",x"18"
		,x"A9",x"1A",x"8D",x"02",x"18",x"4C",x"A7",x"EA"
		,x"AD",x"00",x"18",x"29",x"01",x"D0",x"F9",x"A9"
		,x"01",x"8D",x"05",x"18",x"4C",x"DF",x"E9",x"A9"
		,x"FF",x"85",x"51",x"4C",x"C6",x"C8",x"85",x"FF"
		,x"4C",x"00",x"C1",x"C9",x"02",x"90",x"07",x"C9"
		,x"0F",x"F0",x"03",x"4C",x"6B",x"D3",x"4C",x"73"
		,x"D3",x"78",x"A2",x"45",x"9A",x"4C",x"25",x"EB"
		,x"2C",x"01",x"18",x"4C",x"5B",x"E8",x"BD",x"FF"
		,x"00",x"60",x"A6",x"7F",x"BD",x"FF",x"00",x"4C"
		,x"1B",x"F0",x"A9",x"00",x"9D",x"FF",x"00",x"4C"
		,x"B7",x"C1",x"98",x"9D",x"FF",x"00",x"4C",x"64"
		,x"C6",x"95",x"1C",x"9D",x"FF",x"00",x"4C",x"75"
		,x"D0",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"
		,x"AA",x"AA",x"AA",x"AA",x"AA",x"EB",x"C6",x"C8"
		,x"8F",x"F9",x"5F",x"CD",x"97",x"CD",x"00",x"05"
		,x"03",x"05",x"06",x"05",x"09",x"05",x"0C",x"05"
		,x"0F",x"05",x"01",x"FF",x"A0",x"EA",x"67",x"FE"
			);
begin
	p_rom : process(clk)
	begin
	if clk'event and clk= '0' then
		data <= ROM(to_integer(unsigned(addr)));
	end if;
	end process;
end rtl;
